 // NumberOfConfigBits: 253
module SCC6_switch_matrix
    #(
        parameter NoConfigBits=253
    )
    (
        input i_0to60,
        input i_0to61,
        input i_0to62,
        input i_0to63,
        input i_0to64,
        input i_0to65,
        input i_0to66,
        input i_0to67,
        input i_0to68,
        input i_0to69,
        input i_0to610,
        input i_0to611,
        input i_0to612,
        input i_0to613,
        input i_0to614,
        input i_0to615,
        input i_0to616,
        input i_0to617,
        input i_0to618,
        input i_0to619,
        input i_0to620,
        input i_0to621,
        input i_0to622,
        input i_0to623,
        input i_0to624,
        input i_0to625,
        input i_0to626,
        input i_0to627,
        input i_0to628,
        input i_0to629,
        input i_0to630,
        input i_0to631,
        input i_0to632,
        input i_0to633,
        input i_0to634,
        input i_0to635,
        input i_0to636,
        input i_0to637,
        input i_0to638,
        input i_0to639,
        input i_0to640,
        input i_0to641,
        input i_0to642,
        input i_0to643,
        input i_0to644,
        input i_0to645,
        input i_0to646,
        input i_0to647,
        input i_1to60,
        input i_1to61,
        input i_1to62,
        input i_1to63,
        input i_1to64,
        input i_1to65,
        input i_1to66,
        input i_1to67,
        input i_1to68,
        input i_1to69,
        input i_1to610,
        input i_1to611,
        input i_1to612,
        input i_1to613,
        input i_1to614,
        input i_1to615,
        input i_1to616,
        input i_1to617,
        input i_1to618,
        input i_1to619,
        input i_1to620,
        input i_1to621,
        input i_1to622,
        input i_1to623,
        input i_1to624,
        input i_1to625,
        input i_1to626,
        input i_1to627,
        input i_1to628,
        input i_1to629,
        input i_1to630,
        input i_1to631,
        input i_1to632,
        input i_1to633,
        input i_1to634,
        input i_1to635,
        input i_1to636,
        input i_1to637,
        input i_1to638,
        input i_1to639,
        input i_2to60,
        input i_2to61,
        input i_2to62,
        input i_2to63,
        input i_2to64,
        input i_2to65,
        input i_2to66,
        input i_2to67,
        input i_2to68,
        input i_2to69,
        input i_2to610,
        input i_2to611,
        input i_2to612,
        input i_2to613,
        input i_2to614,
        input i_2to615,
        input i_2to616,
        input i_2to617,
        input i_2to618,
        input i_2to619,
        input i_2to620,
        input i_2to621,
        input i_2to622,
        input i_2to623,
        input i_2to624,
        input i_2to625,
        input i_2to626,
        input i_2to627,
        input i_2to628,
        input i_2to629,
        input i_2to630,
        input i_2to631,
        input i_3to60,
        input i_3to61,
        input i_3to62,
        input i_3to63,
        input i_3to64,
        input i_3to65,
        input i_3to66,
        input i_3to67,
        input i_3to68,
        input i_3to69,
        input i_3to610,
        input i_3to611,
        input i_3to612,
        input i_3to613,
        input i_3to614,
        input i_3to615,
        input i_3to616,
        input i_3to617,
        input i_3to618,
        input i_3to619,
        input i_3to620,
        input i_3to621,
        input i_3to622,
        input i_3to623,
        input i_4to60,
        input i_4to61,
        input i_4to62,
        input i_4to63,
        input i_4to64,
        input i_4to65,
        input i_4to66,
        input i_4to67,
        input i_4to68,
        input i_4to69,
        input i_4to610,
        input i_4to611,
        input i_4to612,
        input i_4to613,
        input i_4to614,
        input i_4to615,
        input i_5to60,
        input i_5to61,
        input i_5to62,
        input i_5to63,
        input i_5to64,
        input i_5to65,
        input i_5to66,
        input i_5to67,
        input i_w2e0,
        input i_w2e1,
        input i_w2e2,
        input i_w2e3,
        input i_w2e4,
        input i_w2e5,
        input i_w2e6,
        input i_w2e7,
        input i_w2e8,
        input i_w2e9,
        input i_w2e10,
        input i_w2e11,
        input i_w2e12,
        input i_w2e13,
        input i_w2e14,
        input i_w2e15,
        input i_w2e16,
        input i_w2e17,
        input i_w2e18,
        input i_w2e19,
        input i_w2e20,
        input i_w2e21,
        input i_w2e22,
        input i_w2e23,
        input i_w2e24,
        input i_w2e25,
        input i_w2e26,
        input i_w2e27,
        input i_w2e28,
        input i_w2e29,
        input i_w2e30,
        input i_w2e31,
        input i_w2e32,
        input i_w2e33,
        input i_w2e34,
        input i_w2e35,
        input i_w2e36,
        input i_w2e37,
        input i_w2e38,
        input i_w2e39,
        input i_w2e40,
        input i_w2e41,
        input i_w2e42,
        input i_w2e43,
        input i_w2e44,
        input i_w2e45,
        input i_w2e46,
        input i_w2e47,
        input i_w2e48,
        input i_w2e49,
        input i_w2e50,
        input i_w2e51,
        input i_w2e52,
        input i_w2e53,
        input i_w2e54,
        input i_w2e55,
        input N1END0,
        input N1END1,
        input N1END2,
        input N1END3,
        input N2MID0,
        input N2MID1,
        input N2MID2,
        input N2MID3,
        input N2MID4,
        input N2MID5,
        input N2MID6,
        input N2MID7,
        input N2END0,
        input N2END1,
        input N2END2,
        input N2END3,
        input N2END4,
        input N2END5,
        input N2END6,
        input N2END7,
        input N4END0,
        input N4END1,
        input N4END2,
        input N4END3,
        input NN4END0,
        input NN4END1,
        input NN4END2,
        input NN4END3,
        input E1END0,
        input E1END1,
        input E1END2,
        input E1END3,
        input E2MID0,
        input E2MID1,
        input E2MID2,
        input E2MID3,
        input E2MID4,
        input E2MID5,
        input E2MID6,
        input E2MID7,
        input E2END0,
        input E2END1,
        input E2END2,
        input E2END3,
        input E2END4,
        input E2END5,
        input E2END6,
        input E2END7,
        input EE4END0,
        input EE4END1,
        input EE4END2,
        input EE4END3,
        input E6END0,
        input E6END1,
        input S1END0,
        input S1END1,
        input S1END2,
        input S1END3,
        input S2MID0,
        input S2MID1,
        input S2MID2,
        input S2MID3,
        input S2MID4,
        input S2MID5,
        input S2MID6,
        input S2MID7,
        input S2END0,
        input S2END1,
        input S2END2,
        input S2END3,
        input S2END4,
        input S2END5,
        input S2END6,
        input S2END7,
        input S4END0,
        input S4END1,
        input S4END2,
        input S4END3,
        input SS4END0,
        input SS4END1,
        input SS4END2,
        input SS4END3,
        input W1END0,
        input W1END1,
        input W1END2,
        input W1END3,
        input W2MID0,
        input W2MID1,
        input W2MID2,
        input W2MID3,
        input W2MID4,
        input W2MID5,
        input W2MID6,
        input W2MID7,
        input W2END0,
        input W2END1,
        input W2END2,
        input W2END3,
        input W2END4,
        input W2END5,
        input W2END6,
        input W2END7,
        input WW4END0,
        input WW4END1,
        input WW4END2,
        input WW4END3,
        input W6END0,
        input W6END1,
        input req_ready,
        input resp_data0,
        input resp_data1,
        input resp_data2,
        input resp_data3,
        input resp_data4,
        input resp_data5,
        input resp_data6,
        input resp_data7,
        input resp_data8,
        input resp_data9,
        input resp_data10,
        input resp_data11,
        input resp_data12,
        input resp_data13,
        input resp_data14,
        input resp_data15,
        input resp_data16,
        input resp_data17,
        input resp_data18,
        input resp_data19,
        input resp_data20,
        input resp_data21,
        input resp_data22,
        input resp_data23,
        input resp_data24,
        input resp_data25,
        input resp_data26,
        input resp_data27,
        input resp_data28,
        input resp_data29,
        input resp_data30,
        input resp_data31,
        input resp_status0,
        input resp_status1,
        input resp_status2,
        input resp_valid,
        input t_req_cxu0,
        input t_req_cxu1,
        input t_req_data00,
        input t_req_data01,
        input t_req_data02,
        input t_req_data03,
        input t_req_data04,
        input t_req_data05,
        input t_req_data06,
        input t_req_data07,
        input t_req_data08,
        input t_req_data09,
        input t_req_data010,
        input t_req_data011,
        input t_req_data012,
        input t_req_data013,
        input t_req_data014,
        input t_req_data015,
        input t_req_data016,
        input t_req_data017,
        input t_req_data018,
        input t_req_data019,
        input t_req_data020,
        input t_req_data021,
        input t_req_data022,
        input t_req_data023,
        input t_req_data024,
        input t_req_data025,
        input t_req_data026,
        input t_req_data027,
        input t_req_data028,
        input t_req_data029,
        input t_req_data030,
        input t_req_data031,
        input t_req_data10,
        input t_req_data11,
        input t_req_data12,
        input t_req_data13,
        input t_req_data14,
        input t_req_data15,
        input t_req_data16,
        input t_req_data17,
        input t_req_data18,
        input t_req_data19,
        input t_req_data110,
        input t_req_data111,
        input t_req_data112,
        input t_req_data113,
        input t_req_data114,
        input t_req_data115,
        input t_req_data116,
        input t_req_data117,
        input t_req_data118,
        input t_req_data119,
        input t_req_data120,
        input t_req_data121,
        input t_req_data122,
        input t_req_data123,
        input t_req_data124,
        input t_req_data125,
        input t_req_data126,
        input t_req_data127,
        input t_req_data128,
        input t_req_data129,
        input t_req_data130,
        input t_req_data131,
        input t_req_func0,
        input t_req_func1,
        input t_req_func2,
        input t_req_insn,
        input t_req_state,
        input t_req_valid,
        input t_resp_ready,
        input J2MID_ABa_END0,
        input J2MID_ABa_END1,
        input J2MID_ABa_END2,
        input J2MID_ABa_END3,
        input J2MID_CDa_END0,
        input J2MID_CDa_END1,
        input J2MID_CDa_END2,
        input J2MID_CDa_END3,
        input J2MID_EFa_END0,
        input J2MID_EFa_END1,
        input J2MID_EFa_END2,
        input J2MID_EFa_END3,
        input J2MID_GHa_END0,
        input J2MID_GHa_END1,
        input J2MID_GHa_END2,
        input J2MID_GHa_END3,
        input J2MID_ABb_END0,
        input J2MID_ABb_END1,
        input J2MID_ABb_END2,
        input J2MID_ABb_END3,
        input J2MID_CDb_END0,
        input J2MID_CDb_END1,
        input J2MID_CDb_END2,
        input J2MID_CDb_END3,
        input J2MID_EFb_END0,
        input J2MID_EFb_END1,
        input J2MID_EFb_END2,
        input J2MID_EFb_END3,
        input J2MID_GHb_END0,
        input J2MID_GHb_END1,
        input J2MID_GHb_END2,
        input J2MID_GHb_END3,
        input J2END_AB_END0,
        input J2END_AB_END1,
        input J2END_AB_END2,
        input J2END_AB_END3,
        input J2END_CD_END0,
        input J2END_CD_END1,
        input J2END_CD_END2,
        input J2END_CD_END3,
        input J2END_EF_END0,
        input J2END_EF_END1,
        input J2END_EF_END2,
        input J2END_EF_END3,
        input J2END_GH_END0,
        input J2END_GH_END1,
        input J2END_GH_END2,
        input J2END_GH_END3,
        input JN2END0,
        input JN2END1,
        input JN2END2,
        input JN2END3,
        input JN2END4,
        input JN2END5,
        input JN2END6,
        input JN2END7,
        input JE2END0,
        input JE2END1,
        input JE2END2,
        input JE2END3,
        input JE2END4,
        input JE2END5,
        input JE2END6,
        input JE2END7,
        input JS2END0,
        input JS2END1,
        input JS2END2,
        input JS2END3,
        input JS2END4,
        input JS2END5,
        input JS2END6,
        input JS2END7,
        input JW2END0,
        input JW2END1,
        input JW2END2,
        input JW2END3,
        input JW2END4,
        input JW2END5,
        input JW2END6,
        input JW2END7,
        input J_l_AB_END0,
        input J_l_AB_END1,
        input J_l_AB_END2,
        input J_l_AB_END3,
        input J_l_CD_END0,
        input J_l_CD_END1,
        input J_l_CD_END2,
        input J_l_CD_END3,
        input J_l_EF_END0,
        input J_l_EF_END1,
        input J_l_EF_END2,
        input J_l_EF_END3,
        input J_l_GH_END0,
        input J_l_GH_END1,
        input J_l_GH_END2,
        input J_l_GH_END3,
        output o_6to00,
        output o_6to01,
        output o_6to02,
        output o_6to03,
        output o_6to04,
        output o_6to05,
        output o_6to06,
        output o_6to07,
        output o_6to08,
        output o_6to09,
        output o_6to010,
        output o_6to011,
        output o_6to012,
        output o_6to013,
        output o_6to014,
        output o_6to015,
        output o_6to016,
        output o_6to017,
        output o_6to018,
        output o_6to019,
        output o_6to020,
        output o_6to021,
        output o_6to022,
        output o_6to023,
        output o_6to024,
        output o_6to025,
        output o_6to026,
        output o_6to027,
        output o_6to028,
        output o_6to029,
        output o_6to030,
        output o_6to031,
        output o_6to032,
        output o_6to033,
        output o_6to034,
        output o_6to035,
        output o_6to036,
        output o_6to037,
        output o_6to038,
        output o_6to039,
        output o_6to040,
        output o_6to041,
        output o_6to042,
        output o_6to043,
        output o_6to044,
        output o_6to045,
        output o_6to046,
        output o_6to047,
        output o_6to10,
        output o_6to11,
        output o_6to12,
        output o_6to13,
        output o_6to14,
        output o_6to15,
        output o_6to16,
        output o_6to17,
        output o_6to18,
        output o_6to19,
        output o_6to110,
        output o_6to111,
        output o_6to112,
        output o_6to113,
        output o_6to114,
        output o_6to115,
        output o_6to116,
        output o_6to117,
        output o_6to118,
        output o_6to119,
        output o_6to120,
        output o_6to121,
        output o_6to122,
        output o_6to123,
        output o_6to124,
        output o_6to125,
        output o_6to126,
        output o_6to127,
        output o_6to128,
        output o_6to129,
        output o_6to130,
        output o_6to131,
        output o_6to132,
        output o_6to133,
        output o_6to134,
        output o_6to135,
        output o_6to136,
        output o_6to137,
        output o_6to138,
        output o_6to139,
        output o_6to20,
        output o_6to21,
        output o_6to22,
        output o_6to23,
        output o_6to24,
        output o_6to25,
        output o_6to26,
        output o_6to27,
        output o_6to28,
        output o_6to29,
        output o_6to210,
        output o_6to211,
        output o_6to212,
        output o_6to213,
        output o_6to214,
        output o_6to215,
        output o_6to216,
        output o_6to217,
        output o_6to218,
        output o_6to219,
        output o_6to220,
        output o_6to221,
        output o_6to222,
        output o_6to223,
        output o_6to224,
        output o_6to225,
        output o_6to226,
        output o_6to227,
        output o_6to228,
        output o_6to229,
        output o_6to230,
        output o_6to231,
        output o_6to30,
        output o_6to31,
        output o_6to32,
        output o_6to33,
        output o_6to34,
        output o_6to35,
        output o_6to36,
        output o_6to37,
        output o_6to38,
        output o_6to39,
        output o_6to310,
        output o_6to311,
        output o_6to312,
        output o_6to313,
        output o_6to314,
        output o_6to315,
        output o_6to316,
        output o_6to317,
        output o_6to318,
        output o_6to319,
        output o_6to320,
        output o_6to321,
        output o_6to322,
        output o_6to323,
        output o_6to40,
        output o_6to41,
        output o_6to42,
        output o_6to43,
        output o_6to44,
        output o_6to45,
        output o_6to46,
        output o_6to47,
        output o_6to48,
        output o_6to49,
        output o_6to410,
        output o_6to411,
        output o_6to412,
        output o_6to413,
        output o_6to414,
        output o_6to415,
        output o_6to50,
        output o_6to51,
        output o_6to52,
        output o_6to53,
        output o_6to54,
        output o_6to55,
        output o_6to56,
        output o_6to57,
        output o_e2w0,
        output o_e2w1,
        output o_e2w2,
        output o_e2w3,
        output o_e2w4,
        output o_e2w5,
        output o_e2w6,
        output o_e2w7,
        output o_e2w8,
        output o_e2w9,
        output o_e2w10,
        output o_e2w11,
        output o_e2w12,
        output o_e2w13,
        output o_e2w14,
        output o_e2w15,
        output o_e2w16,
        output o_e2w17,
        output o_e2w18,
        output o_e2w19,
        output o_e2w20,
        output o_e2w21,
        output o_e2w22,
        output o_e2w23,
        output o_e2w24,
        output o_e2w25,
        output o_e2w26,
        output o_e2w27,
        output o_e2w28,
        output o_e2w29,
        output o_e2w30,
        output o_e2w31,
        output o_e2w32,
        output o_e2w33,
        output o_e2w34,
        output o_e2w35,
        output o_e2w36,
        output o_e2w37,
        output o_e2w38,
        output o_e2w39,
        output o_e2w40,
        output o_e2w41,
        output o_e2w42,
        output o_e2w43,
        output o_e2w44,
        output o_e2w45,
        output o_e2w46,
        output o_e2w47,
        output o_e2w48,
        output o_e2w49,
        output o_e2w50,
        output o_e2w51,
        output o_e2w52,
        output o_e2w53,
        output o_e2w54,
        output o_e2w55,
        output N1BEG0,
        output N1BEG1,
        output N1BEG2,
        output N1BEG3,
        output N2BEG0,
        output N2BEG1,
        output N2BEG2,
        output N2BEG3,
        output N2BEG4,
        output N2BEG5,
        output N2BEG6,
        output N2BEG7,
        output N2BEGb0,
        output N2BEGb1,
        output N2BEGb2,
        output N2BEGb3,
        output N2BEGb4,
        output N2BEGb5,
        output N2BEGb6,
        output N2BEGb7,
        output N4BEG0,
        output N4BEG1,
        output N4BEG2,
        output N4BEG3,
        output NN4BEG0,
        output NN4BEG1,
        output NN4BEG2,
        output NN4BEG3,
        output E1BEG0,
        output E1BEG1,
        output E1BEG2,
        output E1BEG3,
        output E2BEG0,
        output E2BEG1,
        output E2BEG2,
        output E2BEG3,
        output E2BEG4,
        output E2BEG5,
        output E2BEG6,
        output E2BEG7,
        output E2BEGb0,
        output E2BEGb1,
        output E2BEGb2,
        output E2BEGb3,
        output E2BEGb4,
        output E2BEGb5,
        output E2BEGb6,
        output E2BEGb7,
        output EE4BEG0,
        output EE4BEG1,
        output EE4BEG2,
        output EE4BEG3,
        output E6BEG0,
        output E6BEG1,
        output S1BEG0,
        output S1BEG1,
        output S1BEG2,
        output S1BEG3,
        output S2BEG0,
        output S2BEG1,
        output S2BEG2,
        output S2BEG3,
        output S2BEG4,
        output S2BEG5,
        output S2BEG6,
        output S2BEG7,
        output S2BEGb0,
        output S2BEGb1,
        output S2BEGb2,
        output S2BEGb3,
        output S2BEGb4,
        output S2BEGb5,
        output S2BEGb6,
        output S2BEGb7,
        output S4BEG0,
        output S4BEG1,
        output S4BEG2,
        output S4BEG3,
        output SS4BEG0,
        output SS4BEG1,
        output SS4BEG2,
        output SS4BEG3,
        output W1BEG0,
        output W1BEG1,
        output W1BEG2,
        output W1BEG3,
        output W2BEG0,
        output W2BEG1,
        output W2BEG2,
        output W2BEG3,
        output W2BEG4,
        output W2BEG5,
        output W2BEG6,
        output W2BEG7,
        output W2BEGb0,
        output W2BEGb1,
        output W2BEGb2,
        output W2BEGb3,
        output W2BEGb4,
        output W2BEGb5,
        output W2BEGb6,
        output W2BEGb7,
        output WW4BEG0,
        output WW4BEG1,
        output WW4BEG2,
        output WW4BEG3,
        output W6BEG0,
        output W6BEG1,
        output clk,
        output clk_en,
        output req_cxu0,
        output req_cxu1,
        output req_data00,
        output req_data01,
        output req_data02,
        output req_data03,
        output req_data04,
        output req_data05,
        output req_data06,
        output req_data07,
        output req_data08,
        output req_data09,
        output req_data010,
        output req_data011,
        output req_data012,
        output req_data013,
        output req_data014,
        output req_data015,
        output req_data016,
        output req_data017,
        output req_data018,
        output req_data019,
        output req_data020,
        output req_data021,
        output req_data022,
        output req_data023,
        output req_data024,
        output req_data025,
        output req_data026,
        output req_data027,
        output req_data028,
        output req_data029,
        output req_data030,
        output req_data031,
        output req_data10,
        output req_data11,
        output req_data12,
        output req_data13,
        output req_data14,
        output req_data15,
        output req_data16,
        output req_data17,
        output req_data18,
        output req_data19,
        output req_data110,
        output req_data111,
        output req_data112,
        output req_data113,
        output req_data114,
        output req_data115,
        output req_data116,
        output req_data117,
        output req_data118,
        output req_data119,
        output req_data120,
        output req_data121,
        output req_data122,
        output req_data123,
        output req_data124,
        output req_data125,
        output req_data126,
        output req_data127,
        output req_data128,
        output req_data129,
        output req_data130,
        output req_data131,
        output req_func0,
        output req_func1,
        output req_func2,
        output req_insn,
        output req_state,
        output req_valid,
        output resp_ready,
        output rst,
        output t_req_ready,
        output t_resp_data0,
        output t_resp_data1,
        output t_resp_data2,
        output t_resp_data3,
        output t_resp_data4,
        output t_resp_data5,
        output t_resp_data6,
        output t_resp_data7,
        output t_resp_data8,
        output t_resp_data9,
        output t_resp_data10,
        output t_resp_data11,
        output t_resp_data12,
        output t_resp_data13,
        output t_resp_data14,
        output t_resp_data15,
        output t_resp_data16,
        output t_resp_data17,
        output t_resp_data18,
        output t_resp_data19,
        output t_resp_data20,
        output t_resp_data21,
        output t_resp_data22,
        output t_resp_data23,
        output t_resp_data24,
        output t_resp_data25,
        output t_resp_data26,
        output t_resp_data27,
        output t_resp_data28,
        output t_resp_data29,
        output t_resp_data30,
        output t_resp_data31,
        output t_resp_status0,
        output t_resp_status1,
        output t_resp_status2,
        output t_resp_valid,
        output J2MID_ABa_BEG0,
        output J2MID_ABa_BEG1,
        output J2MID_ABa_BEG2,
        output J2MID_ABa_BEG3,
        output J2MID_CDa_BEG0,
        output J2MID_CDa_BEG1,
        output J2MID_CDa_BEG2,
        output J2MID_CDa_BEG3,
        output J2MID_EFa_BEG0,
        output J2MID_EFa_BEG1,
        output J2MID_EFa_BEG2,
        output J2MID_EFa_BEG3,
        output J2MID_GHa_BEG0,
        output J2MID_GHa_BEG1,
        output J2MID_GHa_BEG2,
        output J2MID_GHa_BEG3,
        output J2MID_ABb_BEG0,
        output J2MID_ABb_BEG1,
        output J2MID_ABb_BEG2,
        output J2MID_ABb_BEG3,
        output J2MID_CDb_BEG0,
        output J2MID_CDb_BEG1,
        output J2MID_CDb_BEG2,
        output J2MID_CDb_BEG3,
        output J2MID_EFb_BEG0,
        output J2MID_EFb_BEG1,
        output J2MID_EFb_BEG2,
        output J2MID_EFb_BEG3,
        output J2MID_GHb_BEG0,
        output J2MID_GHb_BEG1,
        output J2MID_GHb_BEG2,
        output J2MID_GHb_BEG3,
        output J2END_AB_BEG0,
        output J2END_AB_BEG1,
        output J2END_AB_BEG2,
        output J2END_AB_BEG3,
        output J2END_CD_BEG0,
        output J2END_CD_BEG1,
        output J2END_CD_BEG2,
        output J2END_CD_BEG3,
        output J2END_EF_BEG0,
        output J2END_EF_BEG1,
        output J2END_EF_BEG2,
        output J2END_EF_BEG3,
        output J2END_GH_BEG0,
        output J2END_GH_BEG1,
        output J2END_GH_BEG2,
        output J2END_GH_BEG3,
        output JN2BEG0,
        output JN2BEG1,
        output JN2BEG2,
        output JN2BEG3,
        output JN2BEG4,
        output JN2BEG5,
        output JN2BEG6,
        output JN2BEG7,
        output JE2BEG0,
        output JE2BEG1,
        output JE2BEG2,
        output JE2BEG3,
        output JE2BEG4,
        output JE2BEG5,
        output JE2BEG6,
        output JE2BEG7,
        output JS2BEG0,
        output JS2BEG1,
        output JS2BEG2,
        output JS2BEG3,
        output JS2BEG4,
        output JS2BEG5,
        output JS2BEG6,
        output JS2BEG7,
        output JW2BEG0,
        output JW2BEG1,
        output JW2BEG2,
        output JW2BEG3,
        output JW2BEG4,
        output JW2BEG5,
        output JW2BEG6,
        output JW2BEG7,
        output J_l_AB_BEG0,
        output J_l_AB_BEG1,
        output J_l_AB_BEG2,
        output J_l_AB_BEG3,
        output J_l_CD_BEG0,
        output J_l_CD_BEG1,
        output J_l_CD_BEG2,
        output J_l_CD_BEG3,
        output J_l_EF_BEG0,
        output J_l_EF_BEG1,
        output J_l_EF_BEG2,
        output J_l_EF_BEG3,
        output J_l_GH_BEG0,
        output J_l_GH_BEG1,
        output J_l_GH_BEG2,
        output J_l_GH_BEG3,
 //global
        input [NoConfigBits-1:0] ConfigBits,
        input [NoConfigBits-1:0] ConfigBits_N
);
parameter GND0 = 1'b0;
parameter GND = 1'b0;
parameter VCC0 = 1'b1;
parameter VCC = 1'b1;
parameter VDD0 = 1'b1;
parameter VDD = 1'b1;

wire[1-1:0] o_6to00_input;
wire[1-1:0] o_6to01_input;
wire[1-1:0] o_6to02_input;
wire[1-1:0] o_6to03_input;
wire[1-1:0] o_6to04_input;
wire[1-1:0] o_6to05_input;
wire[1-1:0] o_6to06_input;
wire[1-1:0] o_6to07_input;
wire[0-1:0] o_6to08_input;
wire[0-1:0] o_6to09_input;
wire[0-1:0] o_6to010_input;
wire[0-1:0] o_6to011_input;
wire[0-1:0] o_6to012_input;
wire[0-1:0] o_6to013_input;
wire[0-1:0] o_6to014_input;
wire[0-1:0] o_6to015_input;
wire[0-1:0] o_6to016_input;
wire[0-1:0] o_6to017_input;
wire[0-1:0] o_6to018_input;
wire[0-1:0] o_6to019_input;
wire[0-1:0] o_6to020_input;
wire[0-1:0] o_6to021_input;
wire[0-1:0] o_6to022_input;
wire[0-1:0] o_6to023_input;
wire[0-1:0] o_6to024_input;
wire[0-1:0] o_6to025_input;
wire[0-1:0] o_6to026_input;
wire[0-1:0] o_6to027_input;
wire[0-1:0] o_6to028_input;
wire[0-1:0] o_6to029_input;
wire[0-1:0] o_6to030_input;
wire[0-1:0] o_6to031_input;
wire[0-1:0] o_6to032_input;
wire[0-1:0] o_6to033_input;
wire[0-1:0] o_6to034_input;
wire[0-1:0] o_6to035_input;
wire[0-1:0] o_6to036_input;
wire[0-1:0] o_6to037_input;
wire[0-1:0] o_6to038_input;
wire[0-1:0] o_6to039_input;
wire[0-1:0] o_6to040_input;
wire[0-1:0] o_6to041_input;
wire[0-1:0] o_6to042_input;
wire[0-1:0] o_6to043_input;
wire[0-1:0] o_6to044_input;
wire[0-1:0] o_6to045_input;
wire[0-1:0] o_6to046_input;
wire[0-1:0] o_6to047_input;
wire[1-1:0] o_6to10_input;
wire[1-1:0] o_6to11_input;
wire[1-1:0] o_6to12_input;
wire[1-1:0] o_6to13_input;
wire[1-1:0] o_6to14_input;
wire[1-1:0] o_6to15_input;
wire[1-1:0] o_6to16_input;
wire[1-1:0] o_6to17_input;
wire[0-1:0] o_6to18_input;
wire[0-1:0] o_6to19_input;
wire[0-1:0] o_6to110_input;
wire[0-1:0] o_6to111_input;
wire[0-1:0] o_6to112_input;
wire[0-1:0] o_6to113_input;
wire[0-1:0] o_6to114_input;
wire[0-1:0] o_6to115_input;
wire[0-1:0] o_6to116_input;
wire[0-1:0] o_6to117_input;
wire[0-1:0] o_6to118_input;
wire[0-1:0] o_6to119_input;
wire[0-1:0] o_6to120_input;
wire[0-1:0] o_6to121_input;
wire[0-1:0] o_6to122_input;
wire[0-1:0] o_6to123_input;
wire[0-1:0] o_6to124_input;
wire[0-1:0] o_6to125_input;
wire[0-1:0] o_6to126_input;
wire[0-1:0] o_6to127_input;
wire[0-1:0] o_6to128_input;
wire[0-1:0] o_6to129_input;
wire[0-1:0] o_6to130_input;
wire[0-1:0] o_6to131_input;
wire[0-1:0] o_6to132_input;
wire[0-1:0] o_6to133_input;
wire[0-1:0] o_6to134_input;
wire[0-1:0] o_6to135_input;
wire[0-1:0] o_6to136_input;
wire[0-1:0] o_6to137_input;
wire[0-1:0] o_6to138_input;
wire[0-1:0] o_6to139_input;
wire[1-1:0] o_6to20_input;
wire[1-1:0] o_6to21_input;
wire[1-1:0] o_6to22_input;
wire[1-1:0] o_6to23_input;
wire[1-1:0] o_6to24_input;
wire[1-1:0] o_6to25_input;
wire[1-1:0] o_6to26_input;
wire[1-1:0] o_6to27_input;
wire[0-1:0] o_6to28_input;
wire[0-1:0] o_6to29_input;
wire[0-1:0] o_6to210_input;
wire[0-1:0] o_6to211_input;
wire[0-1:0] o_6to212_input;
wire[0-1:0] o_6to213_input;
wire[0-1:0] o_6to214_input;
wire[0-1:0] o_6to215_input;
wire[0-1:0] o_6to216_input;
wire[0-1:0] o_6to217_input;
wire[0-1:0] o_6to218_input;
wire[0-1:0] o_6to219_input;
wire[0-1:0] o_6to220_input;
wire[0-1:0] o_6to221_input;
wire[0-1:0] o_6to222_input;
wire[0-1:0] o_6to223_input;
wire[0-1:0] o_6to224_input;
wire[0-1:0] o_6to225_input;
wire[0-1:0] o_6to226_input;
wire[0-1:0] o_6to227_input;
wire[0-1:0] o_6to228_input;
wire[0-1:0] o_6to229_input;
wire[0-1:0] o_6to230_input;
wire[0-1:0] o_6to231_input;
wire[1-1:0] o_6to30_input;
wire[1-1:0] o_6to31_input;
wire[1-1:0] o_6to32_input;
wire[1-1:0] o_6to33_input;
wire[1-1:0] o_6to34_input;
wire[1-1:0] o_6to35_input;
wire[1-1:0] o_6to36_input;
wire[1-1:0] o_6to37_input;
wire[0-1:0] o_6to38_input;
wire[0-1:0] o_6to39_input;
wire[0-1:0] o_6to310_input;
wire[0-1:0] o_6to311_input;
wire[0-1:0] o_6to312_input;
wire[0-1:0] o_6to313_input;
wire[0-1:0] o_6to314_input;
wire[0-1:0] o_6to315_input;
wire[0-1:0] o_6to316_input;
wire[0-1:0] o_6to317_input;
wire[0-1:0] o_6to318_input;
wire[0-1:0] o_6to319_input;
wire[0-1:0] o_6to320_input;
wire[0-1:0] o_6to321_input;
wire[0-1:0] o_6to322_input;
wire[0-1:0] o_6to323_input;
wire[1-1:0] o_6to40_input;
wire[1-1:0] o_6to41_input;
wire[1-1:0] o_6to42_input;
wire[1-1:0] o_6to43_input;
wire[1-1:0] o_6to44_input;
wire[1-1:0] o_6to45_input;
wire[1-1:0] o_6to46_input;
wire[1-1:0] o_6to47_input;
wire[0-1:0] o_6to48_input;
wire[0-1:0] o_6to49_input;
wire[0-1:0] o_6to410_input;
wire[0-1:0] o_6to411_input;
wire[0-1:0] o_6to412_input;
wire[0-1:0] o_6to413_input;
wire[0-1:0] o_6to414_input;
wire[0-1:0] o_6to415_input;
wire[1-1:0] o_6to50_input;
wire[1-1:0] o_6to51_input;
wire[1-1:0] o_6to52_input;
wire[1-1:0] o_6to53_input;
wire[1-1:0] o_6to54_input;
wire[1-1:0] o_6to55_input;
wire[1-1:0] o_6to56_input;
wire[1-1:0] o_6to57_input;
wire[1-1:0] o_e2w0_input;
wire[1-1:0] o_e2w1_input;
wire[1-1:0] o_e2w2_input;
wire[1-1:0] o_e2w3_input;
wire[1-1:0] o_e2w4_input;
wire[1-1:0] o_e2w5_input;
wire[1-1:0] o_e2w6_input;
wire[1-1:0] o_e2w7_input;
wire[1-1:0] o_e2w8_input;
wire[1-1:0] o_e2w9_input;
wire[1-1:0] o_e2w10_input;
wire[1-1:0] o_e2w11_input;
wire[1-1:0] o_e2w12_input;
wire[1-1:0] o_e2w13_input;
wire[1-1:0] o_e2w14_input;
wire[1-1:0] o_e2w15_input;
wire[1-1:0] o_e2w16_input;
wire[1-1:0] o_e2w17_input;
wire[1-1:0] o_e2w18_input;
wire[1-1:0] o_e2w19_input;
wire[1-1:0] o_e2w20_input;
wire[1-1:0] o_e2w21_input;
wire[1-1:0] o_e2w22_input;
wire[1-1:0] o_e2w23_input;
wire[1-1:0] o_e2w24_input;
wire[1-1:0] o_e2w25_input;
wire[1-1:0] o_e2w26_input;
wire[1-1:0] o_e2w27_input;
wire[1-1:0] o_e2w28_input;
wire[1-1:0] o_e2w29_input;
wire[1-1:0] o_e2w30_input;
wire[1-1:0] o_e2w31_input;
wire[1-1:0] o_e2w32_input;
wire[1-1:0] o_e2w33_input;
wire[1-1:0] o_e2w34_input;
wire[1-1:0] o_e2w35_input;
wire[1-1:0] o_e2w36_input;
wire[1-1:0] o_e2w37_input;
wire[1-1:0] o_e2w38_input;
wire[1-1:0] o_e2w39_input;
wire[1-1:0] o_e2w40_input;
wire[1-1:0] o_e2w41_input;
wire[1-1:0] o_e2w42_input;
wire[1-1:0] o_e2w43_input;
wire[1-1:0] o_e2w44_input;
wire[1-1:0] o_e2w45_input;
wire[1-1:0] o_e2w46_input;
wire[1-1:0] o_e2w47_input;
wire[1-1:0] o_e2w48_input;
wire[1-1:0] o_e2w49_input;
wire[1-1:0] o_e2w50_input;
wire[1-1:0] o_e2w51_input;
wire[1-1:0] o_e2w52_input;
wire[1-1:0] o_e2w53_input;
wire[1-1:0] o_e2w54_input;
wire[1-1:0] o_e2w55_input;
wire[4-1:0] N1BEG0_input;
wire[4-1:0] N1BEG1_input;
wire[4-1:0] N1BEG2_input;
wire[4-1:0] N1BEG3_input;
wire[1-1:0] N2BEG0_input;
wire[1-1:0] N2BEG1_input;
wire[1-1:0] N2BEG2_input;
wire[1-1:0] N2BEG3_input;
wire[1-1:0] N2BEG4_input;
wire[1-1:0] N2BEG5_input;
wire[1-1:0] N2BEG6_input;
wire[1-1:0] N2BEG7_input;
wire[1-1:0] N2BEGb0_input;
wire[1-1:0] N2BEGb1_input;
wire[1-1:0] N2BEGb2_input;
wire[1-1:0] N2BEGb3_input;
wire[1-1:0] N2BEGb4_input;
wire[1-1:0] N2BEGb5_input;
wire[1-1:0] N2BEGb6_input;
wire[1-1:0] N2BEGb7_input;
wire[4-1:0] N4BEG0_input;
wire[4-1:0] N4BEG1_input;
wire[4-1:0] N4BEG2_input;
wire[4-1:0] N4BEG3_input;
wire[8-1:0] NN4BEG0_input;
wire[8-1:0] NN4BEG1_input;
wire[8-1:0] NN4BEG2_input;
wire[8-1:0] NN4BEG3_input;
wire[4-1:0] E1BEG0_input;
wire[4-1:0] E1BEG1_input;
wire[4-1:0] E1BEG2_input;
wire[4-1:0] E1BEG3_input;
wire[1-1:0] E2BEG0_input;
wire[1-1:0] E2BEG1_input;
wire[1-1:0] E2BEG2_input;
wire[1-1:0] E2BEG3_input;
wire[1-1:0] E2BEG4_input;
wire[1-1:0] E2BEG5_input;
wire[1-1:0] E2BEG6_input;
wire[1-1:0] E2BEG7_input;
wire[1-1:0] E2BEGb0_input;
wire[1-1:0] E2BEGb1_input;
wire[1-1:0] E2BEGb2_input;
wire[1-1:0] E2BEGb3_input;
wire[1-1:0] E2BEGb4_input;
wire[1-1:0] E2BEGb5_input;
wire[1-1:0] E2BEGb6_input;
wire[1-1:0] E2BEGb7_input;
wire[8-1:0] EE4BEG0_input;
wire[8-1:0] EE4BEG1_input;
wire[8-1:0] EE4BEG2_input;
wire[8-1:0] EE4BEG3_input;
wire[16-1:0] E6BEG0_input;
wire[16-1:0] E6BEG1_input;
wire[4-1:0] S1BEG0_input;
wire[4-1:0] S1BEG1_input;
wire[4-1:0] S1BEG2_input;
wire[4-1:0] S1BEG3_input;
wire[1-1:0] S2BEG0_input;
wire[1-1:0] S2BEG1_input;
wire[1-1:0] S2BEG2_input;
wire[1-1:0] S2BEG3_input;
wire[1-1:0] S2BEG4_input;
wire[1-1:0] S2BEG5_input;
wire[1-1:0] S2BEG6_input;
wire[1-1:0] S2BEG7_input;
wire[1-1:0] S2BEGb0_input;
wire[1-1:0] S2BEGb1_input;
wire[1-1:0] S2BEGb2_input;
wire[1-1:0] S2BEGb3_input;
wire[1-1:0] S2BEGb4_input;
wire[1-1:0] S2BEGb5_input;
wire[1-1:0] S2BEGb6_input;
wire[1-1:0] S2BEGb7_input;
wire[4-1:0] S4BEG0_input;
wire[4-1:0] S4BEG1_input;
wire[4-1:0] S4BEG2_input;
wire[4-1:0] S4BEG3_input;
wire[8-1:0] SS4BEG0_input;
wire[8-1:0] SS4BEG1_input;
wire[8-1:0] SS4BEG2_input;
wire[8-1:0] SS4BEG3_input;
wire[4-1:0] W1BEG0_input;
wire[4-1:0] W1BEG1_input;
wire[4-1:0] W1BEG2_input;
wire[4-1:0] W1BEG3_input;
wire[1-1:0] W2BEG0_input;
wire[1-1:0] W2BEG1_input;
wire[1-1:0] W2BEG2_input;
wire[1-1:0] W2BEG3_input;
wire[1-1:0] W2BEG4_input;
wire[1-1:0] W2BEG5_input;
wire[1-1:0] W2BEG6_input;
wire[1-1:0] W2BEG7_input;
wire[1-1:0] W2BEGb0_input;
wire[1-1:0] W2BEGb1_input;
wire[1-1:0] W2BEGb2_input;
wire[1-1:0] W2BEGb3_input;
wire[1-1:0] W2BEGb4_input;
wire[1-1:0] W2BEGb5_input;
wire[1-1:0] W2BEGb6_input;
wire[1-1:0] W2BEGb7_input;
wire[8-1:0] WW4BEG0_input;
wire[8-1:0] WW4BEG1_input;
wire[8-1:0] WW4BEG2_input;
wire[8-1:0] WW4BEG3_input;
wire[16-1:0] W6BEG0_input;
wire[16-1:0] W6BEG1_input;
wire[0-1:0] clk_input;
wire[0-1:0] clk_en_input;
wire[1-1:0] req_cxu0_input;
wire[1-1:0] req_cxu1_input;
wire[1-1:0] req_data00_input;
wire[1-1:0] req_data01_input;
wire[1-1:0] req_data02_input;
wire[1-1:0] req_data03_input;
wire[1-1:0] req_data04_input;
wire[1-1:0] req_data05_input;
wire[1-1:0] req_data06_input;
wire[1-1:0] req_data07_input;
wire[1-1:0] req_data08_input;
wire[1-1:0] req_data09_input;
wire[1-1:0] req_data010_input;
wire[1-1:0] req_data011_input;
wire[1-1:0] req_data012_input;
wire[1-1:0] req_data013_input;
wire[1-1:0] req_data014_input;
wire[1-1:0] req_data015_input;
wire[1-1:0] req_data016_input;
wire[1-1:0] req_data017_input;
wire[1-1:0] req_data018_input;
wire[1-1:0] req_data019_input;
wire[1-1:0] req_data020_input;
wire[1-1:0] req_data021_input;
wire[1-1:0] req_data022_input;
wire[1-1:0] req_data023_input;
wire[1-1:0] req_data024_input;
wire[1-1:0] req_data025_input;
wire[1-1:0] req_data026_input;
wire[1-1:0] req_data027_input;
wire[1-1:0] req_data028_input;
wire[1-1:0] req_data029_input;
wire[1-1:0] req_data030_input;
wire[1-1:0] req_data031_input;
wire[1-1:0] req_data10_input;
wire[1-1:0] req_data11_input;
wire[1-1:0] req_data12_input;
wire[1-1:0] req_data13_input;
wire[1-1:0] req_data14_input;
wire[1-1:0] req_data15_input;
wire[1-1:0] req_data16_input;
wire[1-1:0] req_data17_input;
wire[1-1:0] req_data18_input;
wire[1-1:0] req_data19_input;
wire[1-1:0] req_data110_input;
wire[1-1:0] req_data111_input;
wire[1-1:0] req_data112_input;
wire[1-1:0] req_data113_input;
wire[1-1:0] req_data114_input;
wire[1-1:0] req_data115_input;
wire[1-1:0] req_data116_input;
wire[1-1:0] req_data117_input;
wire[1-1:0] req_data118_input;
wire[1-1:0] req_data119_input;
wire[1-1:0] req_data120_input;
wire[1-1:0] req_data121_input;
wire[1-1:0] req_data122_input;
wire[1-1:0] req_data123_input;
wire[1-1:0] req_data124_input;
wire[1-1:0] req_data125_input;
wire[1-1:0] req_data126_input;
wire[1-1:0] req_data127_input;
wire[1-1:0] req_data128_input;
wire[1-1:0] req_data129_input;
wire[1-1:0] req_data130_input;
wire[1-1:0] req_data131_input;
wire[1-1:0] req_func0_input;
wire[1-1:0] req_func1_input;
wire[1-1:0] req_func2_input;
wire[1-1:0] req_insn_input;
wire[1-1:0] req_state_input;
wire[1-1:0] req_valid_input;
wire[4-1:0] resp_ready_input;
wire[0-1:0] rst_input;
wire[4-1:0] t_req_ready_input;
wire[1-1:0] t_resp_data0_input;
wire[1-1:0] t_resp_data1_input;
wire[1-1:0] t_resp_data2_input;
wire[1-1:0] t_resp_data3_input;
wire[1-1:0] t_resp_data4_input;
wire[1-1:0] t_resp_data5_input;
wire[1-1:0] t_resp_data6_input;
wire[1-1:0] t_resp_data7_input;
wire[1-1:0] t_resp_data8_input;
wire[1-1:0] t_resp_data9_input;
wire[1-1:0] t_resp_data10_input;
wire[1-1:0] t_resp_data11_input;
wire[1-1:0] t_resp_data12_input;
wire[1-1:0] t_resp_data13_input;
wire[1-1:0] t_resp_data14_input;
wire[1-1:0] t_resp_data15_input;
wire[1-1:0] t_resp_data16_input;
wire[1-1:0] t_resp_data17_input;
wire[1-1:0] t_resp_data18_input;
wire[1-1:0] t_resp_data19_input;
wire[1-1:0] t_resp_data20_input;
wire[1-1:0] t_resp_data21_input;
wire[1-1:0] t_resp_data22_input;
wire[1-1:0] t_resp_data23_input;
wire[1-1:0] t_resp_data24_input;
wire[1-1:0] t_resp_data25_input;
wire[1-1:0] t_resp_data26_input;
wire[1-1:0] t_resp_data27_input;
wire[1-1:0] t_resp_data28_input;
wire[1-1:0] t_resp_data29_input;
wire[1-1:0] t_resp_data30_input;
wire[1-1:0] t_resp_data31_input;
wire[4-1:0] t_resp_status0_input;
wire[4-1:0] t_resp_status1_input;
wire[4-1:0] t_resp_status2_input;
wire[4-1:0] t_resp_valid_input;
wire[4-1:0] J2MID_ABa_BEG0_input;
wire[4-1:0] J2MID_ABa_BEG1_input;
wire[4-1:0] J2MID_ABa_BEG2_input;
wire[4-1:0] J2MID_ABa_BEG3_input;
wire[4-1:0] J2MID_CDa_BEG0_input;
wire[4-1:0] J2MID_CDa_BEG1_input;
wire[4-1:0] J2MID_CDa_BEG2_input;
wire[4-1:0] J2MID_CDa_BEG3_input;
wire[4-1:0] J2MID_EFa_BEG0_input;
wire[4-1:0] J2MID_EFa_BEG1_input;
wire[4-1:0] J2MID_EFa_BEG2_input;
wire[4-1:0] J2MID_EFa_BEG3_input;
wire[4-1:0] J2MID_GHa_BEG0_input;
wire[4-1:0] J2MID_GHa_BEG1_input;
wire[4-1:0] J2MID_GHa_BEG2_input;
wire[4-1:0] J2MID_GHa_BEG3_input;
wire[4-1:0] J2MID_ABb_BEG0_input;
wire[4-1:0] J2MID_ABb_BEG1_input;
wire[4-1:0] J2MID_ABb_BEG2_input;
wire[4-1:0] J2MID_ABb_BEG3_input;
wire[4-1:0] J2MID_CDb_BEG0_input;
wire[4-1:0] J2MID_CDb_BEG1_input;
wire[4-1:0] J2MID_CDb_BEG2_input;
wire[4-1:0] J2MID_CDb_BEG3_input;
wire[4-1:0] J2MID_EFb_BEG0_input;
wire[4-1:0] J2MID_EFb_BEG1_input;
wire[4-1:0] J2MID_EFb_BEG2_input;
wire[4-1:0] J2MID_EFb_BEG3_input;
wire[4-1:0] J2MID_GHb_BEG0_input;
wire[4-1:0] J2MID_GHb_BEG1_input;
wire[4-1:0] J2MID_GHb_BEG2_input;
wire[4-1:0] J2MID_GHb_BEG3_input;
wire[4-1:0] J2END_AB_BEG0_input;
wire[4-1:0] J2END_AB_BEG1_input;
wire[4-1:0] J2END_AB_BEG2_input;
wire[4-1:0] J2END_AB_BEG3_input;
wire[4-1:0] J2END_CD_BEG0_input;
wire[4-1:0] J2END_CD_BEG1_input;
wire[4-1:0] J2END_CD_BEG2_input;
wire[4-1:0] J2END_CD_BEG3_input;
wire[4-1:0] J2END_EF_BEG0_input;
wire[4-1:0] J2END_EF_BEG1_input;
wire[4-1:0] J2END_EF_BEG2_input;
wire[4-1:0] J2END_EF_BEG3_input;
wire[4-1:0] J2END_GH_BEG0_input;
wire[4-1:0] J2END_GH_BEG1_input;
wire[4-1:0] J2END_GH_BEG2_input;
wire[4-1:0] J2END_GH_BEG3_input;
wire[16-1:0] JN2BEG0_input;
wire[16-1:0] JN2BEG1_input;
wire[16-1:0] JN2BEG2_input;
wire[16-1:0] JN2BEG3_input;
wire[16-1:0] JN2BEG4_input;
wire[16-1:0] JN2BEG5_input;
wire[16-1:0] JN2BEG6_input;
wire[16-1:0] JN2BEG7_input;
wire[16-1:0] JE2BEG0_input;
wire[16-1:0] JE2BEG1_input;
wire[16-1:0] JE2BEG2_input;
wire[16-1:0] JE2BEG3_input;
wire[16-1:0] JE2BEG4_input;
wire[16-1:0] JE2BEG5_input;
wire[16-1:0] JE2BEG6_input;
wire[16-1:0] JE2BEG7_input;
wire[15-1:0] JS2BEG0_input;
wire[16-1:0] JS2BEG1_input;
wire[16-1:0] JS2BEG2_input;
wire[15-1:0] JS2BEG3_input;
wire[16-1:0] JS2BEG4_input;
wire[16-1:0] JS2BEG5_input;
wire[16-1:0] JS2BEG6_input;
wire[16-1:0] JS2BEG7_input;
wire[15-1:0] JW2BEG0_input;
wire[16-1:0] JW2BEG1_input;
wire[16-1:0] JW2BEG2_input;
wire[15-1:0] JW2BEG3_input;
wire[16-1:0] JW2BEG4_input;
wire[16-1:0] JW2BEG5_input;
wire[16-1:0] JW2BEG6_input;
wire[16-1:0] JW2BEG7_input;
wire[4-1:0] J_l_AB_BEG0_input;
wire[4-1:0] J_l_AB_BEG1_input;
wire[4-1:0] J_l_AB_BEG2_input;
wire[4-1:0] J_l_AB_BEG3_input;
wire[4-1:0] J_l_CD_BEG0_input;
wire[4-1:0] J_l_CD_BEG1_input;
wire[4-1:0] J_l_CD_BEG2_input;
wire[4-1:0] J_l_CD_BEG3_input;
wire[4-1:0] J_l_EF_BEG0_input;
wire[4-1:0] J_l_EF_BEG1_input;
wire[4-1:0] J_l_EF_BEG2_input;
wire[4-1:0] J_l_EF_BEG3_input;
wire[4-1:0] J_l_GH_BEG0_input;
wire[4-1:0] J_l_GH_BEG1_input;
wire[4-1:0] J_l_GH_BEG2_input;
wire[4-1:0] J_l_GH_BEG3_input;

wire[2-1:0] DEBUG_select_N1BEG0;
wire[2-1:0] DEBUG_select_N1BEG1;
wire[2-1:0] DEBUG_select_N1BEG2;
wire[2-1:0] DEBUG_select_N1BEG3;
wire[2-1:0] DEBUG_select_N4BEG0;
wire[2-1:0] DEBUG_select_N4BEG1;
wire[2-1:0] DEBUG_select_N4BEG2;
wire[2-1:0] DEBUG_select_N4BEG3;
wire[3-1:0] DEBUG_select_NN4BEG0;
wire[3-1:0] DEBUG_select_NN4BEG1;
wire[3-1:0] DEBUG_select_NN4BEG2;
wire[3-1:0] DEBUG_select_NN4BEG3;
wire[2-1:0] DEBUG_select_E1BEG0;
wire[2-1:0] DEBUG_select_E1BEG1;
wire[2-1:0] DEBUG_select_E1BEG2;
wire[2-1:0] DEBUG_select_E1BEG3;
wire[3-1:0] DEBUG_select_EE4BEG0;
wire[3-1:0] DEBUG_select_EE4BEG1;
wire[3-1:0] DEBUG_select_EE4BEG2;
wire[3-1:0] DEBUG_select_EE4BEG3;
wire[4-1:0] DEBUG_select_E6BEG0;
wire[4-1:0] DEBUG_select_E6BEG1;
wire[2-1:0] DEBUG_select_S1BEG0;
wire[2-1:0] DEBUG_select_S1BEG1;
wire[2-1:0] DEBUG_select_S1BEG2;
wire[2-1:0] DEBUG_select_S1BEG3;
wire[2-1:0] DEBUG_select_S4BEG0;
wire[2-1:0] DEBUG_select_S4BEG1;
wire[2-1:0] DEBUG_select_S4BEG2;
wire[2-1:0] DEBUG_select_S4BEG3;
wire[3-1:0] DEBUG_select_SS4BEG0;
wire[3-1:0] DEBUG_select_SS4BEG1;
wire[3-1:0] DEBUG_select_SS4BEG2;
wire[3-1:0] DEBUG_select_SS4BEG3;
wire[2-1:0] DEBUG_select_W1BEG0;
wire[2-1:0] DEBUG_select_W1BEG1;
wire[2-1:0] DEBUG_select_W1BEG2;
wire[2-1:0] DEBUG_select_W1BEG3;
wire[3-1:0] DEBUG_select_WW4BEG0;
wire[3-1:0] DEBUG_select_WW4BEG1;
wire[3-1:0] DEBUG_select_WW4BEG2;
wire[3-1:0] DEBUG_select_WW4BEG3;
wire[4-1:0] DEBUG_select_W6BEG0;
wire[4-1:0] DEBUG_select_W6BEG1;
wire[2-1:0] DEBUG_select_resp_ready;
wire[2-1:0] DEBUG_select_t_req_ready;
wire[2-1:0] DEBUG_select_t_resp_status0;
wire[2-1:0] DEBUG_select_t_resp_status1;
wire[2-1:0] DEBUG_select_t_resp_status2;
wire[2-1:0] DEBUG_select_t_resp_valid;
wire[2-1:0] DEBUG_select_J2MID_ABa_BEG0;
wire[2-1:0] DEBUG_select_J2MID_ABa_BEG1;
wire[2-1:0] DEBUG_select_J2MID_ABa_BEG2;
wire[2-1:0] DEBUG_select_J2MID_ABa_BEG3;
wire[2-1:0] DEBUG_select_J2MID_CDa_BEG0;
wire[2-1:0] DEBUG_select_J2MID_CDa_BEG1;
wire[2-1:0] DEBUG_select_J2MID_CDa_BEG2;
wire[2-1:0] DEBUG_select_J2MID_CDa_BEG3;
wire[2-1:0] DEBUG_select_J2MID_EFa_BEG0;
wire[2-1:0] DEBUG_select_J2MID_EFa_BEG1;
wire[2-1:0] DEBUG_select_J2MID_EFa_BEG2;
wire[2-1:0] DEBUG_select_J2MID_EFa_BEG3;
wire[2-1:0] DEBUG_select_J2MID_GHa_BEG0;
wire[2-1:0] DEBUG_select_J2MID_GHa_BEG1;
wire[2-1:0] DEBUG_select_J2MID_GHa_BEG2;
wire[2-1:0] DEBUG_select_J2MID_GHa_BEG3;
wire[2-1:0] DEBUG_select_J2MID_ABb_BEG0;
wire[2-1:0] DEBUG_select_J2MID_ABb_BEG1;
wire[2-1:0] DEBUG_select_J2MID_ABb_BEG2;
wire[2-1:0] DEBUG_select_J2MID_ABb_BEG3;
wire[2-1:0] DEBUG_select_J2MID_CDb_BEG0;
wire[2-1:0] DEBUG_select_J2MID_CDb_BEG1;
wire[2-1:0] DEBUG_select_J2MID_CDb_BEG2;
wire[2-1:0] DEBUG_select_J2MID_CDb_BEG3;
wire[2-1:0] DEBUG_select_J2MID_EFb_BEG0;
wire[2-1:0] DEBUG_select_J2MID_EFb_BEG1;
wire[2-1:0] DEBUG_select_J2MID_EFb_BEG2;
wire[2-1:0] DEBUG_select_J2MID_EFb_BEG3;
wire[2-1:0] DEBUG_select_J2MID_GHb_BEG0;
wire[2-1:0] DEBUG_select_J2MID_GHb_BEG1;
wire[2-1:0] DEBUG_select_J2MID_GHb_BEG2;
wire[2-1:0] DEBUG_select_J2MID_GHb_BEG3;
wire[2-1:0] DEBUG_select_J2END_AB_BEG0;
wire[2-1:0] DEBUG_select_J2END_AB_BEG1;
wire[2-1:0] DEBUG_select_J2END_AB_BEG2;
wire[2-1:0] DEBUG_select_J2END_AB_BEG3;
wire[2-1:0] DEBUG_select_J2END_CD_BEG0;
wire[2-1:0] DEBUG_select_J2END_CD_BEG1;
wire[2-1:0] DEBUG_select_J2END_CD_BEG2;
wire[2-1:0] DEBUG_select_J2END_CD_BEG3;
wire[2-1:0] DEBUG_select_J2END_EF_BEG0;
wire[2-1:0] DEBUG_select_J2END_EF_BEG1;
wire[2-1:0] DEBUG_select_J2END_EF_BEG2;
wire[2-1:0] DEBUG_select_J2END_EF_BEG3;
wire[2-1:0] DEBUG_select_J2END_GH_BEG0;
wire[2-1:0] DEBUG_select_J2END_GH_BEG1;
wire[2-1:0] DEBUG_select_J2END_GH_BEG2;
wire[2-1:0] DEBUG_select_J2END_GH_BEG3;
wire[4-1:0] DEBUG_select_JN2BEG0;
wire[4-1:0] DEBUG_select_JN2BEG1;
wire[4-1:0] DEBUG_select_JN2BEG2;
wire[4-1:0] DEBUG_select_JN2BEG3;
wire[4-1:0] DEBUG_select_JN2BEG4;
wire[4-1:0] DEBUG_select_JN2BEG5;
wire[4-1:0] DEBUG_select_JN2BEG6;
wire[4-1:0] DEBUG_select_JN2BEG7;
wire[4-1:0] DEBUG_select_JE2BEG0;
wire[4-1:0] DEBUG_select_JE2BEG1;
wire[4-1:0] DEBUG_select_JE2BEG2;
wire[4-1:0] DEBUG_select_JE2BEG3;
wire[4-1:0] DEBUG_select_JE2BEG4;
wire[4-1:0] DEBUG_select_JE2BEG5;
wire[4-1:0] DEBUG_select_JE2BEG6;
wire[4-1:0] DEBUG_select_JE2BEG7;
wire[4-1:0] DEBUG_select_JS2BEG0;
wire[4-1:0] DEBUG_select_JS2BEG1;
wire[4-1:0] DEBUG_select_JS2BEG2;
wire[4-1:0] DEBUG_select_JS2BEG3;
wire[4-1:0] DEBUG_select_JS2BEG4;
wire[4-1:0] DEBUG_select_JS2BEG5;
wire[4-1:0] DEBUG_select_JS2BEG6;
wire[4-1:0] DEBUG_select_JS2BEG7;
wire[4-1:0] DEBUG_select_JW2BEG0;
wire[4-1:0] DEBUG_select_JW2BEG1;
wire[4-1:0] DEBUG_select_JW2BEG2;
wire[4-1:0] DEBUG_select_JW2BEG3;
wire[4-1:0] DEBUG_select_JW2BEG4;
wire[4-1:0] DEBUG_select_JW2BEG5;
wire[4-1:0] DEBUG_select_JW2BEG6;
wire[4-1:0] DEBUG_select_JW2BEG7;
wire[2-1:0] DEBUG_select_J_l_AB_BEG0;
wire[2-1:0] DEBUG_select_J_l_AB_BEG1;
wire[2-1:0] DEBUG_select_J_l_AB_BEG2;
wire[2-1:0] DEBUG_select_J_l_AB_BEG3;
wire[2-1:0] DEBUG_select_J_l_CD_BEG0;
wire[2-1:0] DEBUG_select_J_l_CD_BEG1;
wire[2-1:0] DEBUG_select_J_l_CD_BEG2;
wire[2-1:0] DEBUG_select_J_l_CD_BEG3;
wire[2-1:0] DEBUG_select_J_l_EF_BEG0;
wire[2-1:0] DEBUG_select_J_l_EF_BEG1;
wire[2-1:0] DEBUG_select_J_l_EF_BEG2;
wire[2-1:0] DEBUG_select_J_l_EF_BEG3;
wire[2-1:0] DEBUG_select_J_l_GH_BEG0;
wire[2-1:0] DEBUG_select_J_l_GH_BEG1;
wire[2-1:0] DEBUG_select_J_l_GH_BEG2;
wire[2-1:0] DEBUG_select_J_l_GH_BEG3;
 //The configuration bits (if any) are just a long shift register
 //This shift register is padded to an even number of flops/latches
 //switch matrix multiplexer o_6to00 MUX-1
assign o_6to00 = t_req_data124;

 //switch matrix multiplexer o_6to01 MUX-1
assign o_6to01 = t_req_data125;

 //switch matrix multiplexer o_6to02 MUX-1
assign o_6to02 = t_req_data126;

 //switch matrix multiplexer o_6to03 MUX-1
assign o_6to03 = t_req_data127;

 //switch matrix multiplexer o_6to04 MUX-1
assign o_6to04 = t_req_data128;

 //switch matrix multiplexer o_6to05 MUX-1
assign o_6to05 = t_req_data129;

 //switch matrix multiplexer o_6to06 MUX-1
assign o_6to06 = t_req_data130;

 //switch matrix multiplexer o_6to07 MUX-1
assign o_6to07 = t_req_data131;

 //switch matrix multiplexer o_6to08 MUX-0
 //WARNING unused multiplexer MUX-o_6to08
 //switch matrix multiplexer o_6to09 MUX-0
 //WARNING unused multiplexer MUX-o_6to09
 //switch matrix multiplexer o_6to010 MUX-0
 //WARNING unused multiplexer MUX-o_6to010
 //switch matrix multiplexer o_6to011 MUX-0
 //WARNING unused multiplexer MUX-o_6to011
 //switch matrix multiplexer o_6to012 MUX-0
 //WARNING unused multiplexer MUX-o_6to012
 //switch matrix multiplexer o_6to013 MUX-0
 //WARNING unused multiplexer MUX-o_6to013
 //switch matrix multiplexer o_6to014 MUX-0
 //WARNING unused multiplexer MUX-o_6to014
 //switch matrix multiplexer o_6to015 MUX-0
 //WARNING unused multiplexer MUX-o_6to015
 //switch matrix multiplexer o_6to016 MUX-0
 //WARNING unused multiplexer MUX-o_6to016
 //switch matrix multiplexer o_6to017 MUX-0
 //WARNING unused multiplexer MUX-o_6to017
 //switch matrix multiplexer o_6to018 MUX-0
 //WARNING unused multiplexer MUX-o_6to018
 //switch matrix multiplexer o_6to019 MUX-0
 //WARNING unused multiplexer MUX-o_6to019
 //switch matrix multiplexer o_6to020 MUX-0
 //WARNING unused multiplexer MUX-o_6to020
 //switch matrix multiplexer o_6to021 MUX-0
 //WARNING unused multiplexer MUX-o_6to021
 //switch matrix multiplexer o_6to022 MUX-0
 //WARNING unused multiplexer MUX-o_6to022
 //switch matrix multiplexer o_6to023 MUX-0
 //WARNING unused multiplexer MUX-o_6to023
 //switch matrix multiplexer o_6to024 MUX-0
 //WARNING unused multiplexer MUX-o_6to024
 //switch matrix multiplexer o_6to025 MUX-0
 //WARNING unused multiplexer MUX-o_6to025
 //switch matrix multiplexer o_6to026 MUX-0
 //WARNING unused multiplexer MUX-o_6to026
 //switch matrix multiplexer o_6to027 MUX-0
 //WARNING unused multiplexer MUX-o_6to027
 //switch matrix multiplexer o_6to028 MUX-0
 //WARNING unused multiplexer MUX-o_6to028
 //switch matrix multiplexer o_6to029 MUX-0
 //WARNING unused multiplexer MUX-o_6to029
 //switch matrix multiplexer o_6to030 MUX-0
 //WARNING unused multiplexer MUX-o_6to030
 //switch matrix multiplexer o_6to031 MUX-0
 //WARNING unused multiplexer MUX-o_6to031
 //switch matrix multiplexer o_6to032 MUX-0
 //WARNING unused multiplexer MUX-o_6to032
 //switch matrix multiplexer o_6to033 MUX-0
 //WARNING unused multiplexer MUX-o_6to033
 //switch matrix multiplexer o_6to034 MUX-0
 //WARNING unused multiplexer MUX-o_6to034
 //switch matrix multiplexer o_6to035 MUX-0
 //WARNING unused multiplexer MUX-o_6to035
 //switch matrix multiplexer o_6to036 MUX-0
 //WARNING unused multiplexer MUX-o_6to036
 //switch matrix multiplexer o_6to037 MUX-0
 //WARNING unused multiplexer MUX-o_6to037
 //switch matrix multiplexer o_6to038 MUX-0
 //WARNING unused multiplexer MUX-o_6to038
 //switch matrix multiplexer o_6to039 MUX-0
 //WARNING unused multiplexer MUX-o_6to039
 //switch matrix multiplexer o_6to040 MUX-0
 //WARNING unused multiplexer MUX-o_6to040
 //switch matrix multiplexer o_6to041 MUX-0
 //WARNING unused multiplexer MUX-o_6to041
 //switch matrix multiplexer o_6to042 MUX-0
 //WARNING unused multiplexer MUX-o_6to042
 //switch matrix multiplexer o_6to043 MUX-0
 //WARNING unused multiplexer MUX-o_6to043
 //switch matrix multiplexer o_6to044 MUX-0
 //WARNING unused multiplexer MUX-o_6to044
 //switch matrix multiplexer o_6to045 MUX-0
 //WARNING unused multiplexer MUX-o_6to045
 //switch matrix multiplexer o_6to046 MUX-0
 //WARNING unused multiplexer MUX-o_6to046
 //switch matrix multiplexer o_6to047 MUX-0
 //WARNING unused multiplexer MUX-o_6to047
 //switch matrix multiplexer o_6to10 MUX-1
assign o_6to10 = t_req_data116;

 //switch matrix multiplexer o_6to11 MUX-1
assign o_6to11 = t_req_data117;

 //switch matrix multiplexer o_6to12 MUX-1
assign o_6to12 = t_req_data118;

 //switch matrix multiplexer o_6to13 MUX-1
assign o_6to13 = t_req_data119;

 //switch matrix multiplexer o_6to14 MUX-1
assign o_6to14 = t_req_data120;

 //switch matrix multiplexer o_6to15 MUX-1
assign o_6to15 = t_req_data121;

 //switch matrix multiplexer o_6to16 MUX-1
assign o_6to16 = t_req_data122;

 //switch matrix multiplexer o_6to17 MUX-1
assign o_6to17 = t_req_data123;

 //switch matrix multiplexer o_6to18 MUX-0
 //WARNING unused multiplexer MUX-o_6to18
 //switch matrix multiplexer o_6to19 MUX-0
 //WARNING unused multiplexer MUX-o_6to19
 //switch matrix multiplexer o_6to110 MUX-0
 //WARNING unused multiplexer MUX-o_6to110
 //switch matrix multiplexer o_6to111 MUX-0
 //WARNING unused multiplexer MUX-o_6to111
 //switch matrix multiplexer o_6to112 MUX-0
 //WARNING unused multiplexer MUX-o_6to112
 //switch matrix multiplexer o_6to113 MUX-0
 //WARNING unused multiplexer MUX-o_6to113
 //switch matrix multiplexer o_6to114 MUX-0
 //WARNING unused multiplexer MUX-o_6to114
 //switch matrix multiplexer o_6to115 MUX-0
 //WARNING unused multiplexer MUX-o_6to115
 //switch matrix multiplexer o_6to116 MUX-0
 //WARNING unused multiplexer MUX-o_6to116
 //switch matrix multiplexer o_6to117 MUX-0
 //WARNING unused multiplexer MUX-o_6to117
 //switch matrix multiplexer o_6to118 MUX-0
 //WARNING unused multiplexer MUX-o_6to118
 //switch matrix multiplexer o_6to119 MUX-0
 //WARNING unused multiplexer MUX-o_6to119
 //switch matrix multiplexer o_6to120 MUX-0
 //WARNING unused multiplexer MUX-o_6to120
 //switch matrix multiplexer o_6to121 MUX-0
 //WARNING unused multiplexer MUX-o_6to121
 //switch matrix multiplexer o_6to122 MUX-0
 //WARNING unused multiplexer MUX-o_6to122
 //switch matrix multiplexer o_6to123 MUX-0
 //WARNING unused multiplexer MUX-o_6to123
 //switch matrix multiplexer o_6to124 MUX-0
 //WARNING unused multiplexer MUX-o_6to124
 //switch matrix multiplexer o_6to125 MUX-0
 //WARNING unused multiplexer MUX-o_6to125
 //switch matrix multiplexer o_6to126 MUX-0
 //WARNING unused multiplexer MUX-o_6to126
 //switch matrix multiplexer o_6to127 MUX-0
 //WARNING unused multiplexer MUX-o_6to127
 //switch matrix multiplexer o_6to128 MUX-0
 //WARNING unused multiplexer MUX-o_6to128
 //switch matrix multiplexer o_6to129 MUX-0
 //WARNING unused multiplexer MUX-o_6to129
 //switch matrix multiplexer o_6to130 MUX-0
 //WARNING unused multiplexer MUX-o_6to130
 //switch matrix multiplexer o_6to131 MUX-0
 //WARNING unused multiplexer MUX-o_6to131
 //switch matrix multiplexer o_6to132 MUX-0
 //WARNING unused multiplexer MUX-o_6to132
 //switch matrix multiplexer o_6to133 MUX-0
 //WARNING unused multiplexer MUX-o_6to133
 //switch matrix multiplexer o_6to134 MUX-0
 //WARNING unused multiplexer MUX-o_6to134
 //switch matrix multiplexer o_6to135 MUX-0
 //WARNING unused multiplexer MUX-o_6to135
 //switch matrix multiplexer o_6to136 MUX-0
 //WARNING unused multiplexer MUX-o_6to136
 //switch matrix multiplexer o_6to137 MUX-0
 //WARNING unused multiplexer MUX-o_6to137
 //switch matrix multiplexer o_6to138 MUX-0
 //WARNING unused multiplexer MUX-o_6to138
 //switch matrix multiplexer o_6to139 MUX-0
 //WARNING unused multiplexer MUX-o_6to139
 //switch matrix multiplexer o_6to20 MUX-1
assign o_6to20 = t_req_data18;

 //switch matrix multiplexer o_6to21 MUX-1
assign o_6to21 = t_req_data19;

 //switch matrix multiplexer o_6to22 MUX-1
assign o_6to22 = t_req_data110;

 //switch matrix multiplexer o_6to23 MUX-1
assign o_6to23 = t_req_data111;

 //switch matrix multiplexer o_6to24 MUX-1
assign o_6to24 = t_req_data112;

 //switch matrix multiplexer o_6to25 MUX-1
assign o_6to25 = t_req_data113;

 //switch matrix multiplexer o_6to26 MUX-1
assign o_6to26 = t_req_data114;

 //switch matrix multiplexer o_6to27 MUX-1
assign o_6to27 = t_req_data115;

 //switch matrix multiplexer o_6to28 MUX-0
 //WARNING unused multiplexer MUX-o_6to28
 //switch matrix multiplexer o_6to29 MUX-0
 //WARNING unused multiplexer MUX-o_6to29
 //switch matrix multiplexer o_6to210 MUX-0
 //WARNING unused multiplexer MUX-o_6to210
 //switch matrix multiplexer o_6to211 MUX-0
 //WARNING unused multiplexer MUX-o_6to211
 //switch matrix multiplexer o_6to212 MUX-0
 //WARNING unused multiplexer MUX-o_6to212
 //switch matrix multiplexer o_6to213 MUX-0
 //WARNING unused multiplexer MUX-o_6to213
 //switch matrix multiplexer o_6to214 MUX-0
 //WARNING unused multiplexer MUX-o_6to214
 //switch matrix multiplexer o_6to215 MUX-0
 //WARNING unused multiplexer MUX-o_6to215
 //switch matrix multiplexer o_6to216 MUX-0
 //WARNING unused multiplexer MUX-o_6to216
 //switch matrix multiplexer o_6to217 MUX-0
 //WARNING unused multiplexer MUX-o_6to217
 //switch matrix multiplexer o_6to218 MUX-0
 //WARNING unused multiplexer MUX-o_6to218
 //switch matrix multiplexer o_6to219 MUX-0
 //WARNING unused multiplexer MUX-o_6to219
 //switch matrix multiplexer o_6to220 MUX-0
 //WARNING unused multiplexer MUX-o_6to220
 //switch matrix multiplexer o_6to221 MUX-0
 //WARNING unused multiplexer MUX-o_6to221
 //switch matrix multiplexer o_6to222 MUX-0
 //WARNING unused multiplexer MUX-o_6to222
 //switch matrix multiplexer o_6to223 MUX-0
 //WARNING unused multiplexer MUX-o_6to223
 //switch matrix multiplexer o_6to224 MUX-0
 //WARNING unused multiplexer MUX-o_6to224
 //switch matrix multiplexer o_6to225 MUX-0
 //WARNING unused multiplexer MUX-o_6to225
 //switch matrix multiplexer o_6to226 MUX-0
 //WARNING unused multiplexer MUX-o_6to226
 //switch matrix multiplexer o_6to227 MUX-0
 //WARNING unused multiplexer MUX-o_6to227
 //switch matrix multiplexer o_6to228 MUX-0
 //WARNING unused multiplexer MUX-o_6to228
 //switch matrix multiplexer o_6to229 MUX-0
 //WARNING unused multiplexer MUX-o_6to229
 //switch matrix multiplexer o_6to230 MUX-0
 //WARNING unused multiplexer MUX-o_6to230
 //switch matrix multiplexer o_6to231 MUX-0
 //WARNING unused multiplexer MUX-o_6to231
 //switch matrix multiplexer o_6to30 MUX-1
assign o_6to30 = t_req_data10;

 //switch matrix multiplexer o_6to31 MUX-1
assign o_6to31 = t_req_data11;

 //switch matrix multiplexer o_6to32 MUX-1
assign o_6to32 = t_req_data12;

 //switch matrix multiplexer o_6to33 MUX-1
assign o_6to33 = t_req_data13;

 //switch matrix multiplexer o_6to34 MUX-1
assign o_6to34 = t_req_data14;

 //switch matrix multiplexer o_6to35 MUX-1
assign o_6to35 = t_req_data15;

 //switch matrix multiplexer o_6to36 MUX-1
assign o_6to36 = t_req_data16;

 //switch matrix multiplexer o_6to37 MUX-1
assign o_6to37 = t_req_data17;

 //switch matrix multiplexer o_6to38 MUX-0
 //WARNING unused multiplexer MUX-o_6to38
 //switch matrix multiplexer o_6to39 MUX-0
 //WARNING unused multiplexer MUX-o_6to39
 //switch matrix multiplexer o_6to310 MUX-0
 //WARNING unused multiplexer MUX-o_6to310
 //switch matrix multiplexer o_6to311 MUX-0
 //WARNING unused multiplexer MUX-o_6to311
 //switch matrix multiplexer o_6to312 MUX-0
 //WARNING unused multiplexer MUX-o_6to312
 //switch matrix multiplexer o_6to313 MUX-0
 //WARNING unused multiplexer MUX-o_6to313
 //switch matrix multiplexer o_6to314 MUX-0
 //WARNING unused multiplexer MUX-o_6to314
 //switch matrix multiplexer o_6to315 MUX-0
 //WARNING unused multiplexer MUX-o_6to315
 //switch matrix multiplexer o_6to316 MUX-0
 //WARNING unused multiplexer MUX-o_6to316
 //switch matrix multiplexer o_6to317 MUX-0
 //WARNING unused multiplexer MUX-o_6to317
 //switch matrix multiplexer o_6to318 MUX-0
 //WARNING unused multiplexer MUX-o_6to318
 //switch matrix multiplexer o_6to319 MUX-0
 //WARNING unused multiplexer MUX-o_6to319
 //switch matrix multiplexer o_6to320 MUX-0
 //WARNING unused multiplexer MUX-o_6to320
 //switch matrix multiplexer o_6to321 MUX-0
 //WARNING unused multiplexer MUX-o_6to321
 //switch matrix multiplexer o_6to322 MUX-0
 //WARNING unused multiplexer MUX-o_6to322
 //switch matrix multiplexer o_6to323 MUX-0
 //WARNING unused multiplexer MUX-o_6to323
 //switch matrix multiplexer o_6to40 MUX-1
assign o_6to40 = resp_data8;

 //switch matrix multiplexer o_6to41 MUX-1
assign o_6to41 = resp_data9;

 //switch matrix multiplexer o_6to42 MUX-1
assign o_6to42 = resp_data10;

 //switch matrix multiplexer o_6to43 MUX-1
assign o_6to43 = resp_data11;

 //switch matrix multiplexer o_6to44 MUX-1
assign o_6to44 = resp_data12;

 //switch matrix multiplexer o_6to45 MUX-1
assign o_6to45 = resp_data13;

 //switch matrix multiplexer o_6to46 MUX-1
assign o_6to46 = resp_data14;

 //switch matrix multiplexer o_6to47 MUX-1
assign o_6to47 = resp_data15;

 //switch matrix multiplexer o_6to48 MUX-0
 //WARNING unused multiplexer MUX-o_6to48
 //switch matrix multiplexer o_6to49 MUX-0
 //WARNING unused multiplexer MUX-o_6to49
 //switch matrix multiplexer o_6to410 MUX-0
 //WARNING unused multiplexer MUX-o_6to410
 //switch matrix multiplexer o_6to411 MUX-0
 //WARNING unused multiplexer MUX-o_6to411
 //switch matrix multiplexer o_6to412 MUX-0
 //WARNING unused multiplexer MUX-o_6to412
 //switch matrix multiplexer o_6to413 MUX-0
 //WARNING unused multiplexer MUX-o_6to413
 //switch matrix multiplexer o_6to414 MUX-0
 //WARNING unused multiplexer MUX-o_6to414
 //switch matrix multiplexer o_6to415 MUX-0
 //WARNING unused multiplexer MUX-o_6to415
 //switch matrix multiplexer o_6to50 MUX-1
assign o_6to50 = resp_data0;

 //switch matrix multiplexer o_6to51 MUX-1
assign o_6to51 = resp_data1;

 //switch matrix multiplexer o_6to52 MUX-1
assign o_6to52 = resp_data2;

 //switch matrix multiplexer o_6to53 MUX-1
assign o_6to53 = resp_data3;

 //switch matrix multiplexer o_6to54 MUX-1
assign o_6to54 = resp_data4;

 //switch matrix multiplexer o_6to55 MUX-1
assign o_6to55 = resp_data5;

 //switch matrix multiplexer o_6to56 MUX-1
assign o_6to56 = resp_data6;

 //switch matrix multiplexer o_6to57 MUX-1
assign o_6to57 = resp_data7;

 //switch matrix multiplexer o_e2w0 MUX-1
assign o_e2w0 = t_req_valid;

 //switch matrix multiplexer o_e2w1 MUX-1
assign o_e2w1 = t_req_cxu1;

 //switch matrix multiplexer o_e2w2 MUX-1
assign o_e2w2 = t_req_cxu0;

 //switch matrix multiplexer o_e2w3 MUX-1
assign o_e2w3 = t_req_state;

 //switch matrix multiplexer o_e2w4 MUX-1
assign o_e2w4 = t_req_func2;

 //switch matrix multiplexer o_e2w5 MUX-1
assign o_e2w5 = t_req_func1;

 //switch matrix multiplexer o_e2w6 MUX-1
assign o_e2w6 = t_req_func0;

 //switch matrix multiplexer o_e2w7 MUX-1
assign o_e2w7 = t_req_insn;

 //switch matrix multiplexer o_e2w8 MUX-1
assign o_e2w8 = resp_data8;

 //switch matrix multiplexer o_e2w9 MUX-1
assign o_e2w9 = resp_data9;

 //switch matrix multiplexer o_e2w10 MUX-1
assign o_e2w10 = resp_data10;

 //switch matrix multiplexer o_e2w11 MUX-1
assign o_e2w11 = resp_data11;

 //switch matrix multiplexer o_e2w12 MUX-1
assign o_e2w12 = resp_data12;

 //switch matrix multiplexer o_e2w13 MUX-1
assign o_e2w13 = resp_data13;

 //switch matrix multiplexer o_e2w14 MUX-1
assign o_e2w14 = resp_data14;

 //switch matrix multiplexer o_e2w15 MUX-1
assign o_e2w15 = resp_data15;

 //switch matrix multiplexer o_e2w16 MUX-1
assign o_e2w16 = resp_data24;

 //switch matrix multiplexer o_e2w17 MUX-1
assign o_e2w17 = resp_data25;

 //switch matrix multiplexer o_e2w18 MUX-1
assign o_e2w18 = resp_data26;

 //switch matrix multiplexer o_e2w19 MUX-1
assign o_e2w19 = resp_data27;

 //switch matrix multiplexer o_e2w20 MUX-1
assign o_e2w20 = resp_data28;

 //switch matrix multiplexer o_e2w21 MUX-1
assign o_e2w21 = resp_data29;

 //switch matrix multiplexer o_e2w22 MUX-1
assign o_e2w22 = resp_data30;

 //switch matrix multiplexer o_e2w23 MUX-1
assign o_e2w23 = resp_data31;

 //switch matrix multiplexer o_e2w24 MUX-1
assign o_e2w24 = t_req_data00;

 //switch matrix multiplexer o_e2w25 MUX-1
assign o_e2w25 = t_req_data01;

 //switch matrix multiplexer o_e2w26 MUX-1
assign o_e2w26 = t_req_data02;

 //switch matrix multiplexer o_e2w27 MUX-1
assign o_e2w27 = t_req_data03;

 //switch matrix multiplexer o_e2w28 MUX-1
assign o_e2w28 = t_req_data04;

 //switch matrix multiplexer o_e2w29 MUX-1
assign o_e2w29 = t_req_data05;

 //switch matrix multiplexer o_e2w30 MUX-1
assign o_e2w30 = t_req_data06;

 //switch matrix multiplexer o_e2w31 MUX-1
assign o_e2w31 = t_req_data07;

 //switch matrix multiplexer o_e2w32 MUX-1
assign o_e2w32 = t_req_data08;

 //switch matrix multiplexer o_e2w33 MUX-1
assign o_e2w33 = t_req_data09;

 //switch matrix multiplexer o_e2w34 MUX-1
assign o_e2w34 = t_req_data010;

 //switch matrix multiplexer o_e2w35 MUX-1
assign o_e2w35 = t_req_data011;

 //switch matrix multiplexer o_e2w36 MUX-1
assign o_e2w36 = t_req_data012;

 //switch matrix multiplexer o_e2w37 MUX-1
assign o_e2w37 = t_req_data013;

 //switch matrix multiplexer o_e2w38 MUX-1
assign o_e2w38 = t_req_data014;

 //switch matrix multiplexer o_e2w39 MUX-1
assign o_e2w39 = t_req_data015;

 //switch matrix multiplexer o_e2w40 MUX-1
assign o_e2w40 = t_req_data016;

 //switch matrix multiplexer o_e2w41 MUX-1
assign o_e2w41 = t_req_data017;

 //switch matrix multiplexer o_e2w42 MUX-1
assign o_e2w42 = t_req_data018;

 //switch matrix multiplexer o_e2w43 MUX-1
assign o_e2w43 = t_req_data019;

 //switch matrix multiplexer o_e2w44 MUX-1
assign o_e2w44 = t_req_data020;

 //switch matrix multiplexer o_e2w45 MUX-1
assign o_e2w45 = t_req_data021;

 //switch matrix multiplexer o_e2w46 MUX-1
assign o_e2w46 = t_req_data022;

 //switch matrix multiplexer o_e2w47 MUX-1
assign o_e2w47 = t_req_data023;

 //switch matrix multiplexer o_e2w48 MUX-1
assign o_e2w48 = t_req_data024;

 //switch matrix multiplexer o_e2w49 MUX-1
assign o_e2w49 = t_req_data025;

 //switch matrix multiplexer o_e2w50 MUX-1
assign o_e2w50 = t_req_data026;

 //switch matrix multiplexer o_e2w51 MUX-1
assign o_e2w51 = t_req_data027;

 //switch matrix multiplexer o_e2w52 MUX-1
assign o_e2w52 = t_req_data028;

 //switch matrix multiplexer o_e2w53 MUX-1
assign o_e2w53 = t_req_data029;

 //switch matrix multiplexer o_e2w54 MUX-1
assign o_e2w54 = t_req_data030;

 //switch matrix multiplexer o_e2w55 MUX-1
assign o_e2w55 = t_req_data031;

 //switch matrix multiplexer N1BEG0 MUX-4
assign N1BEG0_input = {J_l_CD_END1,JW2END3,J2MID_CDb_END3,resp_valid};
cus_mux41_buf inst_cus_mux41_buf_N1BEG0 (
    .A0(N1BEG0_input[0]),
    .A1(N1BEG0_input[1]),
    .A2(N1BEG0_input[2]),
    .A3(N1BEG0_input[3]),
    .S0(ConfigBits[0+0]),
    .S0N(ConfigBits_N[0+0]),
    .S1(ConfigBits[0+1]),
    .S1N(ConfigBits_N[0+1]),
    .X(N1BEG0)
);

 //switch matrix multiplexer N1BEG1 MUX-4
assign N1BEG1_input = {J_l_EF_END2,JW2END0,J2MID_EFb_END0,resp_status2};
cus_mux41_buf inst_cus_mux41_buf_N1BEG1 (
    .A0(N1BEG1_input[0]),
    .A1(N1BEG1_input[1]),
    .A2(N1BEG1_input[2]),
    .A3(N1BEG1_input[3]),
    .S0(ConfigBits[2+0]),
    .S0N(ConfigBits_N[2+0]),
    .S1(ConfigBits[2+1]),
    .S1N(ConfigBits_N[2+1]),
    .X(N1BEG1)
);

 //switch matrix multiplexer N1BEG2 MUX-4
assign N1BEG2_input = {J_l_GH_END3,JW2END1,J2MID_GHb_END1,resp_status1};
cus_mux41_buf inst_cus_mux41_buf_N1BEG2 (
    .A0(N1BEG2_input[0]),
    .A1(N1BEG2_input[1]),
    .A2(N1BEG2_input[2]),
    .A3(N1BEG2_input[3]),
    .S0(ConfigBits[4+0]),
    .S0N(ConfigBits_N[4+0]),
    .S1(ConfigBits[4+1]),
    .S1N(ConfigBits_N[4+1]),
    .X(N1BEG2)
);

 //switch matrix multiplexer N1BEG3 MUX-4
assign N1BEG3_input = {J_l_AB_END0,JW2END2,J2MID_ABb_END2,resp_status0};
cus_mux41_buf inst_cus_mux41_buf_N1BEG3 (
    .A0(N1BEG3_input[0]),
    .A1(N1BEG3_input[1]),
    .A2(N1BEG3_input[2]),
    .A3(N1BEG3_input[3]),
    .S0(ConfigBits[6+0]),
    .S0N(ConfigBits_N[6+0]),
    .S1(ConfigBits[6+1]),
    .S1N(ConfigBits_N[6+1]),
    .X(N1BEG3)
);

 //switch matrix multiplexer N2BEG0 MUX-1
assign N2BEG0 = JN2END0;

 //switch matrix multiplexer N2BEG1 MUX-1
assign N2BEG1 = JN2END1;

 //switch matrix multiplexer N2BEG2 MUX-1
assign N2BEG2 = JN2END2;

 //switch matrix multiplexer N2BEG3 MUX-1
assign N2BEG3 = JN2END3;

 //switch matrix multiplexer N2BEG4 MUX-1
assign N2BEG4 = JN2END4;

 //switch matrix multiplexer N2BEG5 MUX-1
assign N2BEG5 = JN2END5;

 //switch matrix multiplexer N2BEG6 MUX-1
assign N2BEG6 = JN2END6;

 //switch matrix multiplexer N2BEG7 MUX-1
assign N2BEG7 = JN2END7;

 //switch matrix multiplexer N2BEGb0 MUX-1
assign N2BEGb0 = N2MID0;

 //switch matrix multiplexer N2BEGb1 MUX-1
assign N2BEGb1 = N2MID1;

 //switch matrix multiplexer N2BEGb2 MUX-1
assign N2BEGb2 = N2MID2;

 //switch matrix multiplexer N2BEGb3 MUX-1
assign N2BEGb3 = N2MID3;

 //switch matrix multiplexer N2BEGb4 MUX-1
assign N2BEGb4 = N2MID4;

 //switch matrix multiplexer N2BEGb5 MUX-1
assign N2BEGb5 = N2MID5;

 //switch matrix multiplexer N2BEGb6 MUX-1
assign N2BEGb6 = N2MID6;

 //switch matrix multiplexer N2BEGb7 MUX-1
assign N2BEGb7 = N2MID7;

 //switch matrix multiplexer N4BEG0 MUX-4
assign N4BEG0_input = {resp_status1,E6END1,N4END1,N2END2};
cus_mux41_buf inst_cus_mux41_buf_N4BEG0 (
    .A0(N4BEG0_input[0]),
    .A1(N4BEG0_input[1]),
    .A2(N4BEG0_input[2]),
    .A3(N4BEG0_input[3]),
    .S0(ConfigBits[8+0]),
    .S0N(ConfigBits_N[8+0]),
    .S1(ConfigBits[8+1]),
    .S1N(ConfigBits_N[8+1]),
    .X(N4BEG0)
);

 //switch matrix multiplexer N4BEG1 MUX-4
assign N4BEG1_input = {resp_status0,E6END0,N4END2,N2END3};
cus_mux41_buf inst_cus_mux41_buf_N4BEG1 (
    .A0(N4BEG1_input[0]),
    .A1(N4BEG1_input[1]),
    .A2(N4BEG1_input[2]),
    .A3(N4BEG1_input[3]),
    .S0(ConfigBits[10+0]),
    .S0N(ConfigBits_N[10+0]),
    .S1(ConfigBits[10+1]),
    .S1N(ConfigBits_N[10+1]),
    .X(N4BEG1)
);

 //switch matrix multiplexer N4BEG2 MUX-4
assign N4BEG2_input = {W6END1,S4END0,N4END3,N2END0};
cus_mux41_buf inst_cus_mux41_buf_N4BEG2 (
    .A0(N4BEG2_input[0]),
    .A1(N4BEG2_input[1]),
    .A2(N4BEG2_input[2]),
    .A3(N4BEG2_input[3]),
    .S0(ConfigBits[12+0]),
    .S0N(ConfigBits_N[12+0]),
    .S1(ConfigBits[12+1]),
    .S1N(ConfigBits_N[12+1]),
    .X(N4BEG2)
);

 //switch matrix multiplexer N4BEG3 MUX-4
assign N4BEG3_input = {W6END0,S4END1,N4END0,N2END1};
cus_mux41_buf inst_cus_mux41_buf_N4BEG3 (
    .A0(N4BEG3_input[0]),
    .A1(N4BEG3_input[1]),
    .A2(N4BEG3_input[2]),
    .A3(N4BEG3_input[3]),
    .S0(ConfigBits[14+0]),
    .S0N(ConfigBits_N[14+0]),
    .S1(ConfigBits[14+1]),
    .S1N(ConfigBits_N[14+1]),
    .X(N4BEG3)
);

 //switch matrix multiplexer NN4BEG0 MUX-8
assign NN4BEG0_input = {J2END_GH_END1,J2MID_CDb_END1,J2MID_ABb_END1,resp_status0,W1END2,S4END0,E1END2,N1END2};
cus_mux81_buf inst_cus_mux81_buf_NN4BEG0 (
    .A0(NN4BEG0_input[0]),
    .A1(NN4BEG0_input[1]),
    .A2(NN4BEG0_input[2]),
    .A3(NN4BEG0_input[3]),
    .A4(NN4BEG0_input[4]),
    .A5(NN4BEG0_input[5]),
    .A6(NN4BEG0_input[6]),
    .A7(NN4BEG0_input[7]),
    .S0(ConfigBits[16+0]),
    .S0N(ConfigBits_N[16+0]),
    .S1(ConfigBits[16+1]),
    .S1N(ConfigBits_N[16+1]),
    .S2(ConfigBits[16+2]),
    .S2N(ConfigBits_N[16+2]),
    .X(NN4BEG0)
);

 //switch matrix multiplexer NN4BEG1 MUX-8
assign NN4BEG1_input = {J2END_EF_END1,J2MID_CDa_END2,J2MID_ABa_END2,t_resp_ready,W1END3,S4END1,E1END3,N1END3};
cus_mux81_buf inst_cus_mux81_buf_NN4BEG1 (
    .A0(NN4BEG1_input[0]),
    .A1(NN4BEG1_input[1]),
    .A2(NN4BEG1_input[2]),
    .A3(NN4BEG1_input[3]),
    .A4(NN4BEG1_input[4]),
    .A5(NN4BEG1_input[5]),
    .A6(NN4BEG1_input[6]),
    .A7(NN4BEG1_input[7]),
    .S0(ConfigBits[19+0]),
    .S0N(ConfigBits_N[19+0]),
    .S1(ConfigBits[19+1]),
    .S1N(ConfigBits_N[19+1]),
    .S2(ConfigBits[19+2]),
    .S2N(ConfigBits_N[19+2]),
    .X(NN4BEG1)
);

 //switch matrix multiplexer NN4BEG2 MUX-8
assign NN4BEG2_input = {J2END_CD_END1,J2MID_GHb_END1,J2MID_EFb_END1,resp_valid,req_ready,W1END0,E1END0,N1END0};
cus_mux81_buf inst_cus_mux81_buf_NN4BEG2 (
    .A0(NN4BEG2_input[0]),
    .A1(NN4BEG2_input[1]),
    .A2(NN4BEG2_input[2]),
    .A3(NN4BEG2_input[3]),
    .A4(NN4BEG2_input[4]),
    .A5(NN4BEG2_input[5]),
    .A6(NN4BEG2_input[6]),
    .A7(NN4BEG2_input[7]),
    .S0(ConfigBits[22+0]),
    .S0N(ConfigBits_N[22+0]),
    .S1(ConfigBits[22+1]),
    .S1N(ConfigBits_N[22+1]),
    .S2(ConfigBits[22+2]),
    .S2N(ConfigBits_N[22+2]),
    .X(NN4BEG2)
);

 //switch matrix multiplexer NN4BEG3 MUX-8
assign NN4BEG3_input = {J2END_AB_END1,J2MID_GHa_END2,J2MID_EFa_END2,resp_status2,resp_status1,W1END1,E1END1,N1END1};
cus_mux81_buf inst_cus_mux81_buf_NN4BEG3 (
    .A0(NN4BEG3_input[0]),
    .A1(NN4BEG3_input[1]),
    .A2(NN4BEG3_input[2]),
    .A3(NN4BEG3_input[3]),
    .A4(NN4BEG3_input[4]),
    .A5(NN4BEG3_input[5]),
    .A6(NN4BEG3_input[6]),
    .A7(NN4BEG3_input[7]),
    .S0(ConfigBits[25+0]),
    .S0N(ConfigBits_N[25+0]),
    .S1(ConfigBits[25+1]),
    .S1N(ConfigBits_N[25+1]),
    .S2(ConfigBits[25+2]),
    .S2N(ConfigBits_N[25+2]),
    .X(NN4BEG3)
);

 //switch matrix multiplexer E1BEG0 MUX-4
assign E1BEG0_input = {J_l_CD_END1,JN2END3,J2MID_CDb_END3,resp_status2};
cus_mux41_buf inst_cus_mux41_buf_E1BEG0 (
    .A0(E1BEG0_input[0]),
    .A1(E1BEG0_input[1]),
    .A2(E1BEG0_input[2]),
    .A3(E1BEG0_input[3]),
    .S0(ConfigBits[28+0]),
    .S0N(ConfigBits_N[28+0]),
    .S1(ConfigBits[28+1]),
    .S1N(ConfigBits_N[28+1]),
    .X(E1BEG0)
);

 //switch matrix multiplexer E1BEG1 MUX-4
assign E1BEG1_input = {J_l_EF_END2,JN2END0,J2MID_EFb_END0,resp_status1};
cus_mux41_buf inst_cus_mux41_buf_E1BEG1 (
    .A0(E1BEG1_input[0]),
    .A1(E1BEG1_input[1]),
    .A2(E1BEG1_input[2]),
    .A3(E1BEG1_input[3]),
    .S0(ConfigBits[30+0]),
    .S0N(ConfigBits_N[30+0]),
    .S1(ConfigBits[30+1]),
    .S1N(ConfigBits_N[30+1]),
    .X(E1BEG1)
);

 //switch matrix multiplexer E1BEG2 MUX-4
assign E1BEG2_input = {J_l_GH_END3,JN2END1,J2MID_GHb_END1,resp_status0};
cus_mux41_buf inst_cus_mux41_buf_E1BEG2 (
    .A0(E1BEG2_input[0]),
    .A1(E1BEG2_input[1]),
    .A2(E1BEG2_input[2]),
    .A3(E1BEG2_input[3]),
    .S0(ConfigBits[32+0]),
    .S0N(ConfigBits_N[32+0]),
    .S1(ConfigBits[32+1]),
    .S1N(ConfigBits_N[32+1]),
    .X(E1BEG2)
);

 //switch matrix multiplexer E1BEG3 MUX-4
assign E1BEG3_input = {J_l_AB_END0,JN2END2,J2MID_ABb_END2,S4END0};
cus_mux41_buf inst_cus_mux41_buf_E1BEG3 (
    .A0(E1BEG3_input[0]),
    .A1(E1BEG3_input[1]),
    .A2(E1BEG3_input[2]),
    .A3(E1BEG3_input[3]),
    .S0(ConfigBits[34+0]),
    .S0N(ConfigBits_N[34+0]),
    .S1(ConfigBits[34+1]),
    .S1N(ConfigBits_N[34+1]),
    .X(E1BEG3)
);

 //switch matrix multiplexer E2BEG0 MUX-1
assign E2BEG0 = JE2END0;

 //switch matrix multiplexer E2BEG1 MUX-1
assign E2BEG1 = JE2END1;

 //switch matrix multiplexer E2BEG2 MUX-1
assign E2BEG2 = JE2END2;

 //switch matrix multiplexer E2BEG3 MUX-1
assign E2BEG3 = JE2END3;

 //switch matrix multiplexer E2BEG4 MUX-1
assign E2BEG4 = JE2END4;

 //switch matrix multiplexer E2BEG5 MUX-1
assign E2BEG5 = JE2END5;

 //switch matrix multiplexer E2BEG6 MUX-1
assign E2BEG6 = JE2END6;

 //switch matrix multiplexer E2BEG7 MUX-1
assign E2BEG7 = JE2END7;

 //switch matrix multiplexer E2BEGb0 MUX-1
assign E2BEGb0 = E2MID0;

 //switch matrix multiplexer E2BEGb1 MUX-1
assign E2BEGb1 = E2MID1;

 //switch matrix multiplexer E2BEGb2 MUX-1
assign E2BEGb2 = E2MID2;

 //switch matrix multiplexer E2BEGb3 MUX-1
assign E2BEGb3 = E2MID3;

 //switch matrix multiplexer E2BEGb4 MUX-1
assign E2BEGb4 = E2MID4;

 //switch matrix multiplexer E2BEGb5 MUX-1
assign E2BEGb5 = E2MID5;

 //switch matrix multiplexer E2BEGb6 MUX-1
assign E2BEGb6 = E2MID6;

 //switch matrix multiplexer E2BEGb7 MUX-1
assign E2BEGb7 = E2MID7;

 //switch matrix multiplexer EE4BEG0 MUX-8
assign EE4BEG0_input = {J2END_GH_END0,J2MID_CDb_END1,J2MID_ABb_END1,resp_status0,S4END0,S1END2,E1END2,N1END2};
cus_mux81_buf inst_cus_mux81_buf_EE4BEG0 (
    .A0(EE4BEG0_input[0]),
    .A1(EE4BEG0_input[1]),
    .A2(EE4BEG0_input[2]),
    .A3(EE4BEG0_input[3]),
    .A4(EE4BEG0_input[4]),
    .A5(EE4BEG0_input[5]),
    .A6(EE4BEG0_input[6]),
    .A7(EE4BEG0_input[7]),
    .S0(ConfigBits[36+0]),
    .S0N(ConfigBits_N[36+0]),
    .S1(ConfigBits[36+1]),
    .S1N(ConfigBits_N[36+1]),
    .S2(ConfigBits[36+2]),
    .S2N(ConfigBits_N[36+2]),
    .X(EE4BEG0)
);

 //switch matrix multiplexer EE4BEG1 MUX-8
assign EE4BEG1_input = {J2END_EF_END0,J2MID_CDa_END2,J2MID_ABa_END2,t_resp_ready,S4END1,S1END3,E1END3,N1END3};
cus_mux81_buf inst_cus_mux81_buf_EE4BEG1 (
    .A0(EE4BEG1_input[0]),
    .A1(EE4BEG1_input[1]),
    .A2(EE4BEG1_input[2]),
    .A3(EE4BEG1_input[3]),
    .A4(EE4BEG1_input[4]),
    .A5(EE4BEG1_input[5]),
    .A6(EE4BEG1_input[6]),
    .A7(EE4BEG1_input[7]),
    .S0(ConfigBits[39+0]),
    .S0N(ConfigBits_N[39+0]),
    .S1(ConfigBits[39+1]),
    .S1N(ConfigBits_N[39+1]),
    .S2(ConfigBits[39+2]),
    .S2N(ConfigBits_N[39+2]),
    .X(EE4BEG1)
);

 //switch matrix multiplexer EE4BEG2 MUX-8
assign EE4BEG2_input = {J2END_CD_END0,J2MID_GHb_END1,J2MID_EFb_END1,resp_valid,req_ready,S1END0,E1END0,N1END0};
cus_mux81_buf inst_cus_mux81_buf_EE4BEG2 (
    .A0(EE4BEG2_input[0]),
    .A1(EE4BEG2_input[1]),
    .A2(EE4BEG2_input[2]),
    .A3(EE4BEG2_input[3]),
    .A4(EE4BEG2_input[4]),
    .A5(EE4BEG2_input[5]),
    .A6(EE4BEG2_input[6]),
    .A7(EE4BEG2_input[7]),
    .S0(ConfigBits[42+0]),
    .S0N(ConfigBits_N[42+0]),
    .S1(ConfigBits[42+1]),
    .S1N(ConfigBits_N[42+1]),
    .S2(ConfigBits[42+2]),
    .S2N(ConfigBits_N[42+2]),
    .X(EE4BEG2)
);

 //switch matrix multiplexer EE4BEG3 MUX-8
assign EE4BEG3_input = {J2END_AB_END0,J2MID_GHa_END2,J2MID_EFa_END2,resp_status2,resp_status1,S1END1,E1END1,N1END1};
cus_mux81_buf inst_cus_mux81_buf_EE4BEG3 (
    .A0(EE4BEG3_input[0]),
    .A1(EE4BEG3_input[1]),
    .A2(EE4BEG3_input[2]),
    .A3(EE4BEG3_input[3]),
    .A4(EE4BEG3_input[4]),
    .A5(EE4BEG3_input[5]),
    .A6(EE4BEG3_input[6]),
    .A7(EE4BEG3_input[7]),
    .S0(ConfigBits[45+0]),
    .S0N(ConfigBits_N[45+0]),
    .S1(ConfigBits[45+1]),
    .S1N(ConfigBits_N[45+1]),
    .S2(ConfigBits[45+2]),
    .S2N(ConfigBits_N[45+2]),
    .X(EE4BEG3)
);

 //switch matrix multiplexer E6BEG0 MUX-16
assign E6BEG0_input = {J2MID_GHb_END1,J2MID_EFb_END1,J2MID_CDb_END1,J2MID_ABb_END1,t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END3,SS4END0,S4END1,S4END0,E1END3,NN4END0};
cus_mux161_buf inst_cus_mux161_buf_E6BEG0 (
    .A0(E6BEG0_input[0]),
    .A1(E6BEG0_input[1]),
    .A2(E6BEG0_input[2]),
    .A3(E6BEG0_input[3]),
    .A4(E6BEG0_input[4]),
    .A5(E6BEG0_input[5]),
    .A6(E6BEG0_input[6]),
    .A7(E6BEG0_input[7]),
    .A8(E6BEG0_input[8]),
    .A9(E6BEG0_input[9]),
    .A10(E6BEG0_input[10]),
    .A11(E6BEG0_input[11]),
    .A12(E6BEG0_input[12]),
    .A13(E6BEG0_input[13]),
    .A14(E6BEG0_input[14]),
    .A15(E6BEG0_input[15]),
    .S0(ConfigBits[48+0]),
    .S0N(ConfigBits_N[48+0]),
    .S1(ConfigBits[48+1]),
    .S1N(ConfigBits_N[48+1]),
    .S2(ConfigBits[48+2]),
    .S2N(ConfigBits_N[48+2]),
    .S3(ConfigBits[48+3]),
    .S3N(ConfigBits_N[48+3]),
    .X(E6BEG0)
);

 //switch matrix multiplexer E6BEG1 MUX-16
assign E6BEG1_input = {J2MID_GHa_END2,J2MID_EFa_END2,J2MID_CDa_END2,J2MID_ABa_END2,t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END2,SS4END3,S4END1,S4END0,E1END2,NN4END3};
cus_mux161_buf inst_cus_mux161_buf_E6BEG1 (
    .A0(E6BEG1_input[0]),
    .A1(E6BEG1_input[1]),
    .A2(E6BEG1_input[2]),
    .A3(E6BEG1_input[3]),
    .A4(E6BEG1_input[4]),
    .A5(E6BEG1_input[5]),
    .A6(E6BEG1_input[6]),
    .A7(E6BEG1_input[7]),
    .A8(E6BEG1_input[8]),
    .A9(E6BEG1_input[9]),
    .A10(E6BEG1_input[10]),
    .A11(E6BEG1_input[11]),
    .A12(E6BEG1_input[12]),
    .A13(E6BEG1_input[13]),
    .A14(E6BEG1_input[14]),
    .A15(E6BEG1_input[15]),
    .S0(ConfigBits[52+0]),
    .S0N(ConfigBits_N[52+0]),
    .S1(ConfigBits[52+1]),
    .S1N(ConfigBits_N[52+1]),
    .S2(ConfigBits[52+2]),
    .S2N(ConfigBits_N[52+2]),
    .S3(ConfigBits[52+3]),
    .S3N(ConfigBits_N[52+3]),
    .X(E6BEG1)
);

 //switch matrix multiplexer S1BEG0 MUX-4
assign S1BEG0_input = {J_l_CD_END1,JE2END3,J2MID_CDb_END3,resp_status1};
cus_mux41_buf inst_cus_mux41_buf_S1BEG0 (
    .A0(S1BEG0_input[0]),
    .A1(S1BEG0_input[1]),
    .A2(S1BEG0_input[2]),
    .A3(S1BEG0_input[3]),
    .S0(ConfigBits[56+0]),
    .S0N(ConfigBits_N[56+0]),
    .S1(ConfigBits[56+1]),
    .S1N(ConfigBits_N[56+1]),
    .X(S1BEG0)
);

 //switch matrix multiplexer S1BEG1 MUX-4
assign S1BEG1_input = {J_l_EF_END2,JE2END0,J2MID_EFb_END0,resp_status0};
cus_mux41_buf inst_cus_mux41_buf_S1BEG1 (
    .A0(S1BEG1_input[0]),
    .A1(S1BEG1_input[1]),
    .A2(S1BEG1_input[2]),
    .A3(S1BEG1_input[3]),
    .S0(ConfigBits[58+0]),
    .S0N(ConfigBits_N[58+0]),
    .S1(ConfigBits[58+1]),
    .S1N(ConfigBits_N[58+1]),
    .X(S1BEG1)
);

 //switch matrix multiplexer S1BEG2 MUX-4
assign S1BEG2_input = {J_l_GH_END3,JE2END1,J2MID_GHb_END1,S4END0};
cus_mux41_buf inst_cus_mux41_buf_S1BEG2 (
    .A0(S1BEG2_input[0]),
    .A1(S1BEG2_input[1]),
    .A2(S1BEG2_input[2]),
    .A3(S1BEG2_input[3]),
    .S0(ConfigBits[60+0]),
    .S0N(ConfigBits_N[60+0]),
    .S1(ConfigBits[60+1]),
    .S1N(ConfigBits_N[60+1]),
    .X(S1BEG2)
);

 //switch matrix multiplexer S1BEG3 MUX-4
assign S1BEG3_input = {J_l_AB_END0,JE2END2,J2MID_ABb_END2,S4END1};
cus_mux41_buf inst_cus_mux41_buf_S1BEG3 (
    .A0(S1BEG3_input[0]),
    .A1(S1BEG3_input[1]),
    .A2(S1BEG3_input[2]),
    .A3(S1BEG3_input[3]),
    .S0(ConfigBits[62+0]),
    .S0N(ConfigBits_N[62+0]),
    .S1(ConfigBits[62+1]),
    .S1N(ConfigBits_N[62+1]),
    .X(S1BEG3)
);

 //switch matrix multiplexer S2BEG0 MUX-1
assign S2BEG0 = JS2END0;

 //switch matrix multiplexer S2BEG1 MUX-1
assign S2BEG1 = JS2END1;

 //switch matrix multiplexer S2BEG2 MUX-1
assign S2BEG2 = JS2END2;

 //switch matrix multiplexer S2BEG3 MUX-1
assign S2BEG3 = JS2END3;

 //switch matrix multiplexer S2BEG4 MUX-1
assign S2BEG4 = JS2END4;

 //switch matrix multiplexer S2BEG5 MUX-1
assign S2BEG5 = JS2END5;

 //switch matrix multiplexer S2BEG6 MUX-1
assign S2BEG6 = JS2END6;

 //switch matrix multiplexer S2BEG7 MUX-1
assign S2BEG7 = JS2END7;

 //switch matrix multiplexer S2BEGb0 MUX-1
assign S2BEGb0 = S2MID0;

 //switch matrix multiplexer S2BEGb1 MUX-1
assign S2BEGb1 = S2MID1;

 //switch matrix multiplexer S2BEGb2 MUX-1
assign S2BEGb2 = S2MID2;

 //switch matrix multiplexer S2BEGb3 MUX-1
assign S2BEGb3 = S2MID3;

 //switch matrix multiplexer S2BEGb4 MUX-1
assign S2BEGb4 = S2MID4;

 //switch matrix multiplexer S2BEGb5 MUX-1
assign S2BEGb5 = S2MID5;

 //switch matrix multiplexer S2BEGb6 MUX-1
assign S2BEGb6 = S2MID6;

 //switch matrix multiplexer S2BEGb7 MUX-1
assign S2BEGb7 = S2MID7;

 //switch matrix multiplexer S4BEG0 MUX-4
assign S4BEG0_input = {t_resp_ready,S4END1,S2END2,E6END1};
cus_mux41_buf inst_cus_mux41_buf_S4BEG0 (
    .A0(S4BEG0_input[0]),
    .A1(S4BEG0_input[1]),
    .A2(S4BEG0_input[2]),
    .A3(S4BEG0_input[3]),
    .S0(ConfigBits[64+0]),
    .S0N(ConfigBits_N[64+0]),
    .S1(ConfigBits[64+1]),
    .S1N(ConfigBits_N[64+1]),
    .X(S4BEG0)
);

 //switch matrix multiplexer S4BEG1 MUX-4
assign S4BEG1_input = {req_ready,S4END2,S2END3,E6END0};
cus_mux41_buf inst_cus_mux41_buf_S4BEG1 (
    .A0(S4BEG1_input[0]),
    .A1(S4BEG1_input[1]),
    .A2(S4BEG1_input[2]),
    .A3(S4BEG1_input[3]),
    .S0(ConfigBits[66+0]),
    .S0N(ConfigBits_N[66+0]),
    .S1(ConfigBits[66+1]),
    .S1N(ConfigBits_N[66+1]),
    .X(S4BEG1)
);

 //switch matrix multiplexer S4BEG2 MUX-4
assign S4BEG2_input = {resp_valid,W6END1,S4END3,S2END0};
cus_mux41_buf inst_cus_mux41_buf_S4BEG2 (
    .A0(S4BEG2_input[0]),
    .A1(S4BEG2_input[1]),
    .A2(S4BEG2_input[2]),
    .A3(S4BEG2_input[3]),
    .S0(ConfigBits[68+0]),
    .S0N(ConfigBits_N[68+0]),
    .S1(ConfigBits[68+1]),
    .S1N(ConfigBits_N[68+1]),
    .X(S4BEG2)
);

 //switch matrix multiplexer S4BEG3 MUX-4
assign S4BEG3_input = {resp_status2,W6END0,S4END0,S2END1};
cus_mux41_buf inst_cus_mux41_buf_S4BEG3 (
    .A0(S4BEG3_input[0]),
    .A1(S4BEG3_input[1]),
    .A2(S4BEG3_input[2]),
    .A3(S4BEG3_input[3]),
    .S0(ConfigBits[70+0]),
    .S0N(ConfigBits_N[70+0]),
    .S1(ConfigBits[70+1]),
    .S1N(ConfigBits_N[70+1]),
    .X(S4BEG3)
);

 //switch matrix multiplexer SS4BEG0 MUX-8
assign SS4BEG0_input = {J2END_GH_END3,J2MID_CDb_END1,J2MID_ABb_END1,resp_status0,W1END2,S4END0,E1END2,N1END2};
cus_mux81_buf inst_cus_mux81_buf_SS4BEG0 (
    .A0(SS4BEG0_input[0]),
    .A1(SS4BEG0_input[1]),
    .A2(SS4BEG0_input[2]),
    .A3(SS4BEG0_input[3]),
    .A4(SS4BEG0_input[4]),
    .A5(SS4BEG0_input[5]),
    .A6(SS4BEG0_input[6]),
    .A7(SS4BEG0_input[7]),
    .S0(ConfigBits[72+0]),
    .S0N(ConfigBits_N[72+0]),
    .S1(ConfigBits[72+1]),
    .S1N(ConfigBits_N[72+1]),
    .S2(ConfigBits[72+2]),
    .S2N(ConfigBits_N[72+2]),
    .X(SS4BEG0)
);

 //switch matrix multiplexer SS4BEG1 MUX-8
assign SS4BEG1_input = {J2END_EF_END3,J2MID_CDa_END2,J2MID_ABa_END2,t_resp_ready,W1END3,S4END1,E1END3,N1END3};
cus_mux81_buf inst_cus_mux81_buf_SS4BEG1 (
    .A0(SS4BEG1_input[0]),
    .A1(SS4BEG1_input[1]),
    .A2(SS4BEG1_input[2]),
    .A3(SS4BEG1_input[3]),
    .A4(SS4BEG1_input[4]),
    .A5(SS4BEG1_input[5]),
    .A6(SS4BEG1_input[6]),
    .A7(SS4BEG1_input[7]),
    .S0(ConfigBits[75+0]),
    .S0N(ConfigBits_N[75+0]),
    .S1(ConfigBits[75+1]),
    .S1N(ConfigBits_N[75+1]),
    .S2(ConfigBits[75+2]),
    .S2N(ConfigBits_N[75+2]),
    .X(SS4BEG1)
);

 //switch matrix multiplexer SS4BEG2 MUX-8
assign SS4BEG2_input = {J2END_CD_END3,J2MID_GHb_END1,J2MID_EFb_END1,resp_valid,req_ready,W1END0,E1END0,N1END0};
cus_mux81_buf inst_cus_mux81_buf_SS4BEG2 (
    .A0(SS4BEG2_input[0]),
    .A1(SS4BEG2_input[1]),
    .A2(SS4BEG2_input[2]),
    .A3(SS4BEG2_input[3]),
    .A4(SS4BEG2_input[4]),
    .A5(SS4BEG2_input[5]),
    .A6(SS4BEG2_input[6]),
    .A7(SS4BEG2_input[7]),
    .S0(ConfigBits[78+0]),
    .S0N(ConfigBits_N[78+0]),
    .S1(ConfigBits[78+1]),
    .S1N(ConfigBits_N[78+1]),
    .S2(ConfigBits[78+2]),
    .S2N(ConfigBits_N[78+2]),
    .X(SS4BEG2)
);

 //switch matrix multiplexer SS4BEG3 MUX-8
assign SS4BEG3_input = {J2END_AB_END3,J2MID_GHa_END2,J2MID_EFa_END2,resp_status2,resp_status1,W1END1,E1END1,N1END1};
cus_mux81_buf inst_cus_mux81_buf_SS4BEG3 (
    .A0(SS4BEG3_input[0]),
    .A1(SS4BEG3_input[1]),
    .A2(SS4BEG3_input[2]),
    .A3(SS4BEG3_input[3]),
    .A4(SS4BEG3_input[4]),
    .A5(SS4BEG3_input[5]),
    .A6(SS4BEG3_input[6]),
    .A7(SS4BEG3_input[7]),
    .S0(ConfigBits[81+0]),
    .S0N(ConfigBits_N[81+0]),
    .S1(ConfigBits[81+1]),
    .S1N(ConfigBits_N[81+1]),
    .S2(ConfigBits[81+2]),
    .S2N(ConfigBits_N[81+2]),
    .X(SS4BEG3)
);

 //switch matrix multiplexer W1BEG0 MUX-4
assign W1BEG0_input = {J_l_CD_END1,JS2END3,J2MID_CDb_END3,resp_status0};
cus_mux41_buf inst_cus_mux41_buf_W1BEG0 (
    .A0(W1BEG0_input[0]),
    .A1(W1BEG0_input[1]),
    .A2(W1BEG0_input[2]),
    .A3(W1BEG0_input[3]),
    .S0(ConfigBits[84+0]),
    .S0N(ConfigBits_N[84+0]),
    .S1(ConfigBits[84+1]),
    .S1N(ConfigBits_N[84+1]),
    .X(W1BEG0)
);

 //switch matrix multiplexer W1BEG1 MUX-4
assign W1BEG1_input = {J_l_EF_END2,JS2END0,J2MID_EFb_END0,S4END0};
cus_mux41_buf inst_cus_mux41_buf_W1BEG1 (
    .A0(W1BEG1_input[0]),
    .A1(W1BEG1_input[1]),
    .A2(W1BEG1_input[2]),
    .A3(W1BEG1_input[3]),
    .S0(ConfigBits[86+0]),
    .S0N(ConfigBits_N[86+0]),
    .S1(ConfigBits[86+1]),
    .S1N(ConfigBits_N[86+1]),
    .X(W1BEG1)
);

 //switch matrix multiplexer W1BEG2 MUX-4
assign W1BEG2_input = {J_l_GH_END3,JS2END1,J2MID_GHb_END1,S4END1};
cus_mux41_buf inst_cus_mux41_buf_W1BEG2 (
    .A0(W1BEG2_input[0]),
    .A1(W1BEG2_input[1]),
    .A2(W1BEG2_input[2]),
    .A3(W1BEG2_input[3]),
    .S0(ConfigBits[88+0]),
    .S0N(ConfigBits_N[88+0]),
    .S1(ConfigBits[88+1]),
    .S1N(ConfigBits_N[88+1]),
    .X(W1BEG2)
);

 //switch matrix multiplexer W1BEG3 MUX-4
assign W1BEG3_input = {J_l_AB_END0,JS2END2,J2MID_ABb_END2,t_resp_ready};
cus_mux41_buf inst_cus_mux41_buf_W1BEG3 (
    .A0(W1BEG3_input[0]),
    .A1(W1BEG3_input[1]),
    .A2(W1BEG3_input[2]),
    .A3(W1BEG3_input[3]),
    .S0(ConfigBits[90+0]),
    .S0N(ConfigBits_N[90+0]),
    .S1(ConfigBits[90+1]),
    .S1N(ConfigBits_N[90+1]),
    .X(W1BEG3)
);

 //switch matrix multiplexer W2BEG0 MUX-1
assign W2BEG0 = JW2END0;

 //switch matrix multiplexer W2BEG1 MUX-1
assign W2BEG1 = JW2END1;

 //switch matrix multiplexer W2BEG2 MUX-1
assign W2BEG2 = JW2END2;

 //switch matrix multiplexer W2BEG3 MUX-1
assign W2BEG3 = JW2END3;

 //switch matrix multiplexer W2BEG4 MUX-1
assign W2BEG4 = JW2END4;

 //switch matrix multiplexer W2BEG5 MUX-1
assign W2BEG5 = JW2END5;

 //switch matrix multiplexer W2BEG6 MUX-1
assign W2BEG6 = JW2END6;

 //switch matrix multiplexer W2BEG7 MUX-1
assign W2BEG7 = JW2END7;

 //switch matrix multiplexer W2BEGb0 MUX-1
assign W2BEGb0 = W2MID0;

 //switch matrix multiplexer W2BEGb1 MUX-1
assign W2BEGb1 = W2MID1;

 //switch matrix multiplexer W2BEGb2 MUX-1
assign W2BEGb2 = W2MID2;

 //switch matrix multiplexer W2BEGb3 MUX-1
assign W2BEGb3 = W2MID3;

 //switch matrix multiplexer W2BEGb4 MUX-1
assign W2BEGb4 = W2MID4;

 //switch matrix multiplexer W2BEGb5 MUX-1
assign W2BEGb5 = W2MID5;

 //switch matrix multiplexer W2BEGb6 MUX-1
assign W2BEGb6 = W2MID6;

 //switch matrix multiplexer W2BEGb7 MUX-1
assign W2BEGb7 = W2MID7;

 //switch matrix multiplexer WW4BEG0 MUX-8
assign WW4BEG0_input = {J2END_GH_END2,J2MID_CDb_END1,J2MID_ABb_END1,resp_status0,W1END2,S4END0,S1END2,N1END2};
cus_mux81_buf inst_cus_mux81_buf_WW4BEG0 (
    .A0(WW4BEG0_input[0]),
    .A1(WW4BEG0_input[1]),
    .A2(WW4BEG0_input[2]),
    .A3(WW4BEG0_input[3]),
    .A4(WW4BEG0_input[4]),
    .A5(WW4BEG0_input[5]),
    .A6(WW4BEG0_input[6]),
    .A7(WW4BEG0_input[7]),
    .S0(ConfigBits[92+0]),
    .S0N(ConfigBits_N[92+0]),
    .S1(ConfigBits[92+1]),
    .S1N(ConfigBits_N[92+1]),
    .S2(ConfigBits[92+2]),
    .S2N(ConfigBits_N[92+2]),
    .X(WW4BEG0)
);

 //switch matrix multiplexer WW4BEG1 MUX-8
assign WW4BEG1_input = {J2END_EF_END2,J2MID_CDa_END2,J2MID_ABa_END2,t_resp_ready,W1END3,S4END1,S1END3,N1END3};
cus_mux81_buf inst_cus_mux81_buf_WW4BEG1 (
    .A0(WW4BEG1_input[0]),
    .A1(WW4BEG1_input[1]),
    .A2(WW4BEG1_input[2]),
    .A3(WW4BEG1_input[3]),
    .A4(WW4BEG1_input[4]),
    .A5(WW4BEG1_input[5]),
    .A6(WW4BEG1_input[6]),
    .A7(WW4BEG1_input[7]),
    .S0(ConfigBits[95+0]),
    .S0N(ConfigBits_N[95+0]),
    .S1(ConfigBits[95+1]),
    .S1N(ConfigBits_N[95+1]),
    .S2(ConfigBits[95+2]),
    .S2N(ConfigBits_N[95+2]),
    .X(WW4BEG1)
);

 //switch matrix multiplexer WW4BEG2 MUX-8
assign WW4BEG2_input = {J2END_CD_END2,J2MID_GHb_END1,J2MID_EFb_END1,resp_valid,req_ready,W1END0,S1END0,N1END0};
cus_mux81_buf inst_cus_mux81_buf_WW4BEG2 (
    .A0(WW4BEG2_input[0]),
    .A1(WW4BEG2_input[1]),
    .A2(WW4BEG2_input[2]),
    .A3(WW4BEG2_input[3]),
    .A4(WW4BEG2_input[4]),
    .A5(WW4BEG2_input[5]),
    .A6(WW4BEG2_input[6]),
    .A7(WW4BEG2_input[7]),
    .S0(ConfigBits[98+0]),
    .S0N(ConfigBits_N[98+0]),
    .S1(ConfigBits[98+1]),
    .S1N(ConfigBits_N[98+1]),
    .S2(ConfigBits[98+2]),
    .S2N(ConfigBits_N[98+2]),
    .X(WW4BEG2)
);

 //switch matrix multiplexer WW4BEG3 MUX-8
assign WW4BEG3_input = {J2END_AB_END2,J2MID_GHa_END2,J2MID_EFa_END2,resp_status2,resp_status1,W1END1,S1END1,N1END1};
cus_mux81_buf inst_cus_mux81_buf_WW4BEG3 (
    .A0(WW4BEG3_input[0]),
    .A1(WW4BEG3_input[1]),
    .A2(WW4BEG3_input[2]),
    .A3(WW4BEG3_input[3]),
    .A4(WW4BEG3_input[4]),
    .A5(WW4BEG3_input[5]),
    .A6(WW4BEG3_input[6]),
    .A7(WW4BEG3_input[7]),
    .S0(ConfigBits[101+0]),
    .S0N(ConfigBits_N[101+0]),
    .S1(ConfigBits[101+1]),
    .S1N(ConfigBits_N[101+1]),
    .S2(ConfigBits[101+2]),
    .S2N(ConfigBits_N[101+2]),
    .X(WW4BEG3)
);

 //switch matrix multiplexer W6BEG0 MUX-16
assign W6BEG0_input = {J2MID_GHb_END1,J2MID_EFb_END1,J2MID_CDb_END1,J2MID_ABb_END1,t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END3,SS4END1,S4END1,S4END0,E1END3,NN4END1};
cus_mux161_buf inst_cus_mux161_buf_W6BEG0 (
    .A0(W6BEG0_input[0]),
    .A1(W6BEG0_input[1]),
    .A2(W6BEG0_input[2]),
    .A3(W6BEG0_input[3]),
    .A4(W6BEG0_input[4]),
    .A5(W6BEG0_input[5]),
    .A6(W6BEG0_input[6]),
    .A7(W6BEG0_input[7]),
    .A8(W6BEG0_input[8]),
    .A9(W6BEG0_input[9]),
    .A10(W6BEG0_input[10]),
    .A11(W6BEG0_input[11]),
    .A12(W6BEG0_input[12]),
    .A13(W6BEG0_input[13]),
    .A14(W6BEG0_input[14]),
    .A15(W6BEG0_input[15]),
    .S0(ConfigBits[104+0]),
    .S0N(ConfigBits_N[104+0]),
    .S1(ConfigBits[104+1]),
    .S1N(ConfigBits_N[104+1]),
    .S2(ConfigBits[104+2]),
    .S2N(ConfigBits_N[104+2]),
    .S3(ConfigBits[104+3]),
    .S3N(ConfigBits_N[104+3]),
    .X(W6BEG0)
);

 //switch matrix multiplexer W6BEG1 MUX-16
assign W6BEG1_input = {J2MID_GHa_END2,J2MID_EFa_END2,J2MID_CDa_END2,J2MID_ABa_END2,t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END2,SS4END2,S4END1,S4END0,E1END2,NN4END2};
cus_mux161_buf inst_cus_mux161_buf_W6BEG1 (
    .A0(W6BEG1_input[0]),
    .A1(W6BEG1_input[1]),
    .A2(W6BEG1_input[2]),
    .A3(W6BEG1_input[3]),
    .A4(W6BEG1_input[4]),
    .A5(W6BEG1_input[5]),
    .A6(W6BEG1_input[6]),
    .A7(W6BEG1_input[7]),
    .A8(W6BEG1_input[8]),
    .A9(W6BEG1_input[9]),
    .A10(W6BEG1_input[10]),
    .A11(W6BEG1_input[11]),
    .A12(W6BEG1_input[12]),
    .A13(W6BEG1_input[13]),
    .A14(W6BEG1_input[14]),
    .A15(W6BEG1_input[15]),
    .S0(ConfigBits[108+0]),
    .S0N(ConfigBits_N[108+0]),
    .S1(ConfigBits[108+1]),
    .S1N(ConfigBits_N[108+1]),
    .S2(ConfigBits[108+2]),
    .S2N(ConfigBits_N[108+2]),
    .S3(ConfigBits[108+3]),
    .S3N(ConfigBits_N[108+3]),
    .X(W6BEG1)
);

 //switch matrix multiplexer clk MUX-0
 //WARNING unused multiplexer MUX-clk
 //switch matrix multiplexer clk_en MUX-0
 //WARNING unused multiplexer MUX-clk_en
 //switch matrix multiplexer req_cxu0 MUX-1
assign req_cxu0 = i_w2e2;

 //switch matrix multiplexer req_cxu1 MUX-1
assign req_cxu1 = i_w2e1;

 //switch matrix multiplexer req_data00 MUX-1
assign req_data00 = i_w2e24;

 //switch matrix multiplexer req_data01 MUX-1
assign req_data01 = i_w2e25;

 //switch matrix multiplexer req_data02 MUX-1
assign req_data02 = i_w2e26;

 //switch matrix multiplexer req_data03 MUX-1
assign req_data03 = i_w2e27;

 //switch matrix multiplexer req_data04 MUX-1
assign req_data04 = i_w2e28;

 //switch matrix multiplexer req_data05 MUX-1
assign req_data05 = i_w2e29;

 //switch matrix multiplexer req_data06 MUX-1
assign req_data06 = i_w2e30;

 //switch matrix multiplexer req_data07 MUX-1
assign req_data07 = i_w2e31;

 //switch matrix multiplexer req_data08 MUX-1
assign req_data08 = i_w2e32;

 //switch matrix multiplexer req_data09 MUX-1
assign req_data09 = i_w2e33;

 //switch matrix multiplexer req_data010 MUX-1
assign req_data010 = i_w2e34;

 //switch matrix multiplexer req_data011 MUX-1
assign req_data011 = i_w2e35;

 //switch matrix multiplexer req_data012 MUX-1
assign req_data012 = i_w2e36;

 //switch matrix multiplexer req_data013 MUX-1
assign req_data013 = i_w2e37;

 //switch matrix multiplexer req_data014 MUX-1
assign req_data014 = i_w2e38;

 //switch matrix multiplexer req_data015 MUX-1
assign req_data015 = i_w2e39;

 //switch matrix multiplexer req_data016 MUX-1
assign req_data016 = i_w2e40;

 //switch matrix multiplexer req_data017 MUX-1
assign req_data017 = i_w2e41;

 //switch matrix multiplexer req_data018 MUX-1
assign req_data018 = i_w2e42;

 //switch matrix multiplexer req_data019 MUX-1
assign req_data019 = i_w2e43;

 //switch matrix multiplexer req_data020 MUX-1
assign req_data020 = i_w2e44;

 //switch matrix multiplexer req_data021 MUX-1
assign req_data021 = i_w2e45;

 //switch matrix multiplexer req_data022 MUX-1
assign req_data022 = i_w2e46;

 //switch matrix multiplexer req_data023 MUX-1
assign req_data023 = i_w2e47;

 //switch matrix multiplexer req_data024 MUX-1
assign req_data024 = i_w2e48;

 //switch matrix multiplexer req_data025 MUX-1
assign req_data025 = i_w2e49;

 //switch matrix multiplexer req_data026 MUX-1
assign req_data026 = i_w2e50;

 //switch matrix multiplexer req_data027 MUX-1
assign req_data027 = i_w2e51;

 //switch matrix multiplexer req_data028 MUX-1
assign req_data028 = i_w2e52;

 //switch matrix multiplexer req_data029 MUX-1
assign req_data029 = i_w2e53;

 //switch matrix multiplexer req_data030 MUX-1
assign req_data030 = i_w2e54;

 //switch matrix multiplexer req_data031 MUX-1
assign req_data031 = i_w2e55;

 //switch matrix multiplexer req_data10 MUX-1
assign req_data10 = i_3to60;

 //switch matrix multiplexer req_data11 MUX-1
assign req_data11 = i_3to61;

 //switch matrix multiplexer req_data12 MUX-1
assign req_data12 = i_3to62;

 //switch matrix multiplexer req_data13 MUX-1
assign req_data13 = i_3to63;

 //switch matrix multiplexer req_data14 MUX-1
assign req_data14 = i_3to64;

 //switch matrix multiplexer req_data15 MUX-1
assign req_data15 = i_3to65;

 //switch matrix multiplexer req_data16 MUX-1
assign req_data16 = i_3to66;

 //switch matrix multiplexer req_data17 MUX-1
assign req_data17 = i_3to67;

 //switch matrix multiplexer req_data18 MUX-1
assign req_data18 = i_2to60;

 //switch matrix multiplexer req_data19 MUX-1
assign req_data19 = i_2to61;

 //switch matrix multiplexer req_data110 MUX-1
assign req_data110 = i_2to62;

 //switch matrix multiplexer req_data111 MUX-1
assign req_data111 = i_2to63;

 //switch matrix multiplexer req_data112 MUX-1
assign req_data112 = i_2to64;

 //switch matrix multiplexer req_data113 MUX-1
assign req_data113 = i_2to65;

 //switch matrix multiplexer req_data114 MUX-1
assign req_data114 = i_2to66;

 //switch matrix multiplexer req_data115 MUX-1
assign req_data115 = i_2to67;

 //switch matrix multiplexer req_data116 MUX-1
assign req_data116 = i_1to60;

 //switch matrix multiplexer req_data117 MUX-1
assign req_data117 = i_1to61;

 //switch matrix multiplexer req_data118 MUX-1
assign req_data118 = i_1to62;

 //switch matrix multiplexer req_data119 MUX-1
assign req_data119 = i_1to63;

 //switch matrix multiplexer req_data120 MUX-1
assign req_data120 = i_1to64;

 //switch matrix multiplexer req_data121 MUX-1
assign req_data121 = i_1to65;

 //switch matrix multiplexer req_data122 MUX-1
assign req_data122 = i_1to66;

 //switch matrix multiplexer req_data123 MUX-1
assign req_data123 = i_1to67;

 //switch matrix multiplexer req_data124 MUX-1
assign req_data124 = i_0to60;

 //switch matrix multiplexer req_data125 MUX-1
assign req_data125 = i_0to61;

 //switch matrix multiplexer req_data126 MUX-1
assign req_data126 = i_0to62;

 //switch matrix multiplexer req_data127 MUX-1
assign req_data127 = i_0to63;

 //switch matrix multiplexer req_data128 MUX-1
assign req_data128 = i_0to64;

 //switch matrix multiplexer req_data129 MUX-1
assign req_data129 = i_0to65;

 //switch matrix multiplexer req_data130 MUX-1
assign req_data130 = i_0to66;

 //switch matrix multiplexer req_data131 MUX-1
assign req_data131 = i_0to67;

 //switch matrix multiplexer req_func0 MUX-1
assign req_func0 = i_w2e6;

 //switch matrix multiplexer req_func1 MUX-1
assign req_func1 = i_w2e5;

 //switch matrix multiplexer req_func2 MUX-1
assign req_func2 = i_w2e4;

 //switch matrix multiplexer req_insn MUX-1
assign req_insn = i_w2e7;

 //switch matrix multiplexer req_state MUX-1
assign req_state = i_w2e3;

 //switch matrix multiplexer req_valid MUX-1
assign req_valid = i_w2e0;

 //switch matrix multiplexer resp_ready MUX-4
assign resp_ready_input = {J_l_AB_END0,J2END_AB_END0,J2MID_ABb_END0,J2MID_ABa_END0};
cus_mux41_buf inst_cus_mux41_buf_resp_ready (
    .A0(resp_ready_input[0]),
    .A1(resp_ready_input[1]),
    .A2(resp_ready_input[2]),
    .A3(resp_ready_input[3]),
    .S0(ConfigBits[112+0]),
    .S0N(ConfigBits_N[112+0]),
    .S1(ConfigBits[112+1]),
    .S1N(ConfigBits_N[112+1]),
    .X(resp_ready)
);

 //switch matrix multiplexer rst MUX-0
 //WARNING unused multiplexer MUX-rst
 //switch matrix multiplexer t_req_ready MUX-4
assign t_req_ready_input = {J_l_AB_END1,J2END_AB_END1,J2MID_ABb_END1,J2MID_ABa_END1};
cus_mux41_buf inst_cus_mux41_buf_t_req_ready (
    .A0(t_req_ready_input[0]),
    .A1(t_req_ready_input[1]),
    .A2(t_req_ready_input[2]),
    .A3(t_req_ready_input[3]),
    .S0(ConfigBits[114+0]),
    .S0N(ConfigBits_N[114+0]),
    .S1(ConfigBits[114+1]),
    .S1N(ConfigBits_N[114+1]),
    .X(t_req_ready)
);

 //switch matrix multiplexer t_resp_data0 MUX-1
assign t_resp_data0 = i_5to60;

 //switch matrix multiplexer t_resp_data1 MUX-1
assign t_resp_data1 = i_5to61;

 //switch matrix multiplexer t_resp_data2 MUX-1
assign t_resp_data2 = i_5to62;

 //switch matrix multiplexer t_resp_data3 MUX-1
assign t_resp_data3 = i_5to63;

 //switch matrix multiplexer t_resp_data4 MUX-1
assign t_resp_data4 = i_5to64;

 //switch matrix multiplexer t_resp_data5 MUX-1
assign t_resp_data5 = i_5to65;

 //switch matrix multiplexer t_resp_data6 MUX-1
assign t_resp_data6 = i_5to66;

 //switch matrix multiplexer t_resp_data7 MUX-1
assign t_resp_data7 = i_5to67;

 //switch matrix multiplexer t_resp_data8 MUX-1
assign t_resp_data8 = i_w2e8;

 //switch matrix multiplexer t_resp_data9 MUX-1
assign t_resp_data9 = i_w2e9;

 //switch matrix multiplexer t_resp_data10 MUX-1
assign t_resp_data10 = i_w2e10;

 //switch matrix multiplexer t_resp_data11 MUX-1
assign t_resp_data11 = i_w2e11;

 //switch matrix multiplexer t_resp_data12 MUX-1
assign t_resp_data12 = i_w2e12;

 //switch matrix multiplexer t_resp_data13 MUX-1
assign t_resp_data13 = i_w2e13;

 //switch matrix multiplexer t_resp_data14 MUX-1
assign t_resp_data14 = i_w2e14;

 //switch matrix multiplexer t_resp_data15 MUX-1
assign t_resp_data15 = i_w2e15;

 //switch matrix multiplexer t_resp_data16 MUX-1
assign t_resp_data16 = i_4to60;

 //switch matrix multiplexer t_resp_data17 MUX-1
assign t_resp_data17 = i_4to61;

 //switch matrix multiplexer t_resp_data18 MUX-1
assign t_resp_data18 = i_4to62;

 //switch matrix multiplexer t_resp_data19 MUX-1
assign t_resp_data19 = i_4to63;

 //switch matrix multiplexer t_resp_data20 MUX-1
assign t_resp_data20 = i_4to64;

 //switch matrix multiplexer t_resp_data21 MUX-1
assign t_resp_data21 = i_4to65;

 //switch matrix multiplexer t_resp_data22 MUX-1
assign t_resp_data22 = i_4to66;

 //switch matrix multiplexer t_resp_data23 MUX-1
assign t_resp_data23 = i_4to67;

 //switch matrix multiplexer t_resp_data24 MUX-1
assign t_resp_data24 = i_w2e16;

 //switch matrix multiplexer t_resp_data25 MUX-1
assign t_resp_data25 = i_w2e17;

 //switch matrix multiplexer t_resp_data26 MUX-1
assign t_resp_data26 = i_w2e18;

 //switch matrix multiplexer t_resp_data27 MUX-1
assign t_resp_data27 = i_w2e19;

 //switch matrix multiplexer t_resp_data28 MUX-1
assign t_resp_data28 = i_w2e20;

 //switch matrix multiplexer t_resp_data29 MUX-1
assign t_resp_data29 = i_w2e21;

 //switch matrix multiplexer t_resp_data30 MUX-1
assign t_resp_data30 = i_w2e22;

 //switch matrix multiplexer t_resp_data31 MUX-1
assign t_resp_data31 = i_w2e23;

 //switch matrix multiplexer t_resp_status0 MUX-4
assign t_resp_status0_input = {J_l_EF_END0,J2END_EF_END0,J2MID_EFb_END0,J2MID_EFa_END0};
cus_mux41_buf inst_cus_mux41_buf_t_resp_status0 (
    .A0(t_resp_status0_input[0]),
    .A1(t_resp_status0_input[1]),
    .A2(t_resp_status0_input[2]),
    .A3(t_resp_status0_input[3]),
    .S0(ConfigBits[116+0]),
    .S0N(ConfigBits_N[116+0]),
    .S1(ConfigBits[116+1]),
    .S1N(ConfigBits_N[116+1]),
    .X(t_resp_status0)
);

 //switch matrix multiplexer t_resp_status1 MUX-4
assign t_resp_status1_input = {J_l_EF_END0,J2END_EF_END0,J2MID_EFb_END0,J2MID_EFa_END0};
cus_mux41_buf inst_cus_mux41_buf_t_resp_status1 (
    .A0(t_resp_status1_input[0]),
    .A1(t_resp_status1_input[1]),
    .A2(t_resp_status1_input[2]),
    .A3(t_resp_status1_input[3]),
    .S0(ConfigBits[118+0]),
    .S0N(ConfigBits_N[118+0]),
    .S1(ConfigBits[118+1]),
    .S1N(ConfigBits_N[118+1]),
    .X(t_resp_status1)
);

 //switch matrix multiplexer t_resp_status2 MUX-4
assign t_resp_status2_input = {J_l_CD_END3,J2END_CD_END3,J2MID_CDb_END3,J2MID_CDa_END3};
cus_mux41_buf inst_cus_mux41_buf_t_resp_status2 (
    .A0(t_resp_status2_input[0]),
    .A1(t_resp_status2_input[1]),
    .A2(t_resp_status2_input[2]),
    .A3(t_resp_status2_input[3]),
    .S0(ConfigBits[120+0]),
    .S0N(ConfigBits_N[120+0]),
    .S1(ConfigBits[120+1]),
    .S1N(ConfigBits_N[120+1]),
    .X(t_resp_status2)
);

 //switch matrix multiplexer t_resp_valid MUX-4
assign t_resp_valid_input = {J_l_CD_END2,J2END_CD_END2,J2MID_CDb_END2,J2MID_CDa_END2};
cus_mux41_buf inst_cus_mux41_buf_t_resp_valid (
    .A0(t_resp_valid_input[0]),
    .A1(t_resp_valid_input[1]),
    .A2(t_resp_valid_input[2]),
    .A3(t_resp_valid_input[3]),
    .S0(ConfigBits[122+0]),
    .S0N(ConfigBits_N[122+0]),
    .S1(ConfigBits[122+1]),
    .S1N(ConfigBits_N[122+1]),
    .X(t_resp_valid)
);

 //switch matrix multiplexer J2MID_ABa_BEG0 MUX-4
assign J2MID_ABa_BEG0_input = {JN2END3,W2MID6,S2MID6,N2MID6};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG0 (
    .A0(J2MID_ABa_BEG0_input[0]),
    .A1(J2MID_ABa_BEG0_input[1]),
    .A2(J2MID_ABa_BEG0_input[2]),
    .A3(J2MID_ABa_BEG0_input[3]),
    .S0(ConfigBits[124+0]),
    .S0N(ConfigBits_N[124+0]),
    .S1(ConfigBits[124+1]),
    .S1N(ConfigBits_N[124+1]),
    .X(J2MID_ABa_BEG0)
);

 //switch matrix multiplexer J2MID_ABa_BEG1 MUX-4
assign J2MID_ABa_BEG1_input = {JE2END3,W2MID2,S2MID2,E2MID2};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG1 (
    .A0(J2MID_ABa_BEG1_input[0]),
    .A1(J2MID_ABa_BEG1_input[1]),
    .A2(J2MID_ABa_BEG1_input[2]),
    .A3(J2MID_ABa_BEG1_input[3]),
    .S0(ConfigBits[126+0]),
    .S0N(ConfigBits_N[126+0]),
    .S1(ConfigBits[126+1]),
    .S1N(ConfigBits_N[126+1]),
    .X(J2MID_ABa_BEG1)
);

 //switch matrix multiplexer J2MID_ABa_BEG2 MUX-4
assign J2MID_ABa_BEG2_input = {JS2END3,W2MID4,E2MID4,N2MID4};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG2 (
    .A0(J2MID_ABa_BEG2_input[0]),
    .A1(J2MID_ABa_BEG2_input[1]),
    .A2(J2MID_ABa_BEG2_input[2]),
    .A3(J2MID_ABa_BEG2_input[3]),
    .S0(ConfigBits[128+0]),
    .S0N(ConfigBits_N[128+0]),
    .S1(ConfigBits[128+1]),
    .S1N(ConfigBits_N[128+1]),
    .X(J2MID_ABa_BEG2)
);

 //switch matrix multiplexer J2MID_ABa_BEG3 MUX-4
assign J2MID_ABa_BEG3_input = {JW2END3,S2MID0,E2MID0,N2MID0};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG3 (
    .A0(J2MID_ABa_BEG3_input[0]),
    .A1(J2MID_ABa_BEG3_input[1]),
    .A2(J2MID_ABa_BEG3_input[2]),
    .A3(J2MID_ABa_BEG3_input[3]),
    .S0(ConfigBits[130+0]),
    .S0N(ConfigBits_N[130+0]),
    .S1(ConfigBits[130+1]),
    .S1N(ConfigBits_N[130+1]),
    .X(J2MID_ABa_BEG3)
);

 //switch matrix multiplexer J2MID_CDa_BEG0 MUX-4
assign J2MID_CDa_BEG0_input = {JN2END4,W2MID6,S2MID6,E2MID6};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG0 (
    .A0(J2MID_CDa_BEG0_input[0]),
    .A1(J2MID_CDa_BEG0_input[1]),
    .A2(J2MID_CDa_BEG0_input[2]),
    .A3(J2MID_CDa_BEG0_input[3]),
    .S0(ConfigBits[132+0]),
    .S0N(ConfigBits_N[132+0]),
    .S1(ConfigBits[132+1]),
    .S1N(ConfigBits_N[132+1]),
    .X(J2MID_CDa_BEG0)
);

 //switch matrix multiplexer J2MID_CDa_BEG1 MUX-4
assign J2MID_CDa_BEG1_input = {JE2END4,W2MID2,E2MID2,N2MID2};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG1 (
    .A0(J2MID_CDa_BEG1_input[0]),
    .A1(J2MID_CDa_BEG1_input[1]),
    .A2(J2MID_CDa_BEG1_input[2]),
    .A3(J2MID_CDa_BEG1_input[3]),
    .S0(ConfigBits[134+0]),
    .S0N(ConfigBits_N[134+0]),
    .S1(ConfigBits[134+1]),
    .S1N(ConfigBits_N[134+1]),
    .X(J2MID_CDa_BEG1)
);

 //switch matrix multiplexer J2MID_CDa_BEG2 MUX-4
assign J2MID_CDa_BEG2_input = {JS2END4,S2MID4,E2MID4,N2MID4};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG2 (
    .A0(J2MID_CDa_BEG2_input[0]),
    .A1(J2MID_CDa_BEG2_input[1]),
    .A2(J2MID_CDa_BEG2_input[2]),
    .A3(J2MID_CDa_BEG2_input[3]),
    .S0(ConfigBits[136+0]),
    .S0N(ConfigBits_N[136+0]),
    .S1(ConfigBits[136+1]),
    .S1N(ConfigBits_N[136+1]),
    .X(J2MID_CDa_BEG2)
);

 //switch matrix multiplexer J2MID_CDa_BEG3 MUX-4
assign J2MID_CDa_BEG3_input = {JW2END4,W2MID0,S2MID0,N2MID0};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG3 (
    .A0(J2MID_CDa_BEG3_input[0]),
    .A1(J2MID_CDa_BEG3_input[1]),
    .A2(J2MID_CDa_BEG3_input[2]),
    .A3(J2MID_CDa_BEG3_input[3]),
    .S0(ConfigBits[138+0]),
    .S0N(ConfigBits_N[138+0]),
    .S1(ConfigBits[138+1]),
    .S1N(ConfigBits_N[138+1]),
    .X(J2MID_CDa_BEG3)
);

 //switch matrix multiplexer J2MID_EFa_BEG0 MUX-4
assign J2MID_EFa_BEG0_input = {JN2END5,W2MID6,E2MID6,N2MID6};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG0 (
    .A0(J2MID_EFa_BEG0_input[0]),
    .A1(J2MID_EFa_BEG0_input[1]),
    .A2(J2MID_EFa_BEG0_input[2]),
    .A3(J2MID_EFa_BEG0_input[3]),
    .S0(ConfigBits[140+0]),
    .S0N(ConfigBits_N[140+0]),
    .S1(ConfigBits[140+1]),
    .S1N(ConfigBits_N[140+1]),
    .X(J2MID_EFa_BEG0)
);

 //switch matrix multiplexer J2MID_EFa_BEG1 MUX-4
assign J2MID_EFa_BEG1_input = {JE2END5,S2MID2,E2MID2,N2MID2};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG1 (
    .A0(J2MID_EFa_BEG1_input[0]),
    .A1(J2MID_EFa_BEG1_input[1]),
    .A2(J2MID_EFa_BEG1_input[2]),
    .A3(J2MID_EFa_BEG1_input[3]),
    .S0(ConfigBits[142+0]),
    .S0N(ConfigBits_N[142+0]),
    .S1(ConfigBits[142+1]),
    .S1N(ConfigBits_N[142+1]),
    .X(J2MID_EFa_BEG1)
);

 //switch matrix multiplexer J2MID_EFa_BEG2 MUX-4
assign J2MID_EFa_BEG2_input = {JS2END5,W2MID4,S2MID4,N2MID4};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG2 (
    .A0(J2MID_EFa_BEG2_input[0]),
    .A1(J2MID_EFa_BEG2_input[1]),
    .A2(J2MID_EFa_BEG2_input[2]),
    .A3(J2MID_EFa_BEG2_input[3]),
    .S0(ConfigBits[144+0]),
    .S0N(ConfigBits_N[144+0]),
    .S1(ConfigBits[144+1]),
    .S1N(ConfigBits_N[144+1]),
    .X(J2MID_EFa_BEG2)
);

 //switch matrix multiplexer J2MID_EFa_BEG3 MUX-4
assign J2MID_EFa_BEG3_input = {JW2END5,W2MID0,S2MID0,E2MID0};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG3 (
    .A0(J2MID_EFa_BEG3_input[0]),
    .A1(J2MID_EFa_BEG3_input[1]),
    .A2(J2MID_EFa_BEG3_input[2]),
    .A3(J2MID_EFa_BEG3_input[3]),
    .S0(ConfigBits[146+0]),
    .S0N(ConfigBits_N[146+0]),
    .S1(ConfigBits[146+1]),
    .S1N(ConfigBits_N[146+1]),
    .X(J2MID_EFa_BEG3)
);

 //switch matrix multiplexer J2MID_GHa_BEG0 MUX-4
assign J2MID_GHa_BEG0_input = {JN2END6,S2MID6,E2MID6,N2MID6};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG0 (
    .A0(J2MID_GHa_BEG0_input[0]),
    .A1(J2MID_GHa_BEG0_input[1]),
    .A2(J2MID_GHa_BEG0_input[2]),
    .A3(J2MID_GHa_BEG0_input[3]),
    .S0(ConfigBits[148+0]),
    .S0N(ConfigBits_N[148+0]),
    .S1(ConfigBits[148+1]),
    .S1N(ConfigBits_N[148+1]),
    .X(J2MID_GHa_BEG0)
);

 //switch matrix multiplexer J2MID_GHa_BEG1 MUX-4
assign J2MID_GHa_BEG1_input = {JE2END6,W2MID2,S2MID2,N2MID2};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG1 (
    .A0(J2MID_GHa_BEG1_input[0]),
    .A1(J2MID_GHa_BEG1_input[1]),
    .A2(J2MID_GHa_BEG1_input[2]),
    .A3(J2MID_GHa_BEG1_input[3]),
    .S0(ConfigBits[150+0]),
    .S0N(ConfigBits_N[150+0]),
    .S1(ConfigBits[150+1]),
    .S1N(ConfigBits_N[150+1]),
    .X(J2MID_GHa_BEG1)
);

 //switch matrix multiplexer J2MID_GHa_BEG2 MUX-4
assign J2MID_GHa_BEG2_input = {JS2END6,W2MID4,S2MID4,E2MID4};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG2 (
    .A0(J2MID_GHa_BEG2_input[0]),
    .A1(J2MID_GHa_BEG2_input[1]),
    .A2(J2MID_GHa_BEG2_input[2]),
    .A3(J2MID_GHa_BEG2_input[3]),
    .S0(ConfigBits[152+0]),
    .S0N(ConfigBits_N[152+0]),
    .S1(ConfigBits[152+1]),
    .S1N(ConfigBits_N[152+1]),
    .X(J2MID_GHa_BEG2)
);

 //switch matrix multiplexer J2MID_GHa_BEG3 MUX-4
assign J2MID_GHa_BEG3_input = {JW2END6,W2MID0,E2MID0,N2MID0};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG3 (
    .A0(J2MID_GHa_BEG3_input[0]),
    .A1(J2MID_GHa_BEG3_input[1]),
    .A2(J2MID_GHa_BEG3_input[2]),
    .A3(J2MID_GHa_BEG3_input[3]),
    .S0(ConfigBits[154+0]),
    .S0N(ConfigBits_N[154+0]),
    .S1(ConfigBits[154+1]),
    .S1N(ConfigBits_N[154+1]),
    .X(J2MID_GHa_BEG3)
);

 //switch matrix multiplexer J2MID_ABb_BEG0 MUX-4
assign J2MID_ABb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG0 (
    .A0(J2MID_ABb_BEG0_input[0]),
    .A1(J2MID_ABb_BEG0_input[1]),
    .A2(J2MID_ABb_BEG0_input[2]),
    .A3(J2MID_ABb_BEG0_input[3]),
    .S0(ConfigBits[156+0]),
    .S0N(ConfigBits_N[156+0]),
    .S1(ConfigBits[156+1]),
    .S1N(ConfigBits_N[156+1]),
    .X(J2MID_ABb_BEG0)
);

 //switch matrix multiplexer J2MID_ABb_BEG1 MUX-4
assign J2MID_ABb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG1 (
    .A0(J2MID_ABb_BEG1_input[0]),
    .A1(J2MID_ABb_BEG1_input[1]),
    .A2(J2MID_ABb_BEG1_input[2]),
    .A3(J2MID_ABb_BEG1_input[3]),
    .S0(ConfigBits[158+0]),
    .S0N(ConfigBits_N[158+0]),
    .S1(ConfigBits[158+1]),
    .S1N(ConfigBits_N[158+1]),
    .X(J2MID_ABb_BEG1)
);

 //switch matrix multiplexer J2MID_ABb_BEG2 MUX-4
assign J2MID_ABb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG2 (
    .A0(J2MID_ABb_BEG2_input[0]),
    .A1(J2MID_ABb_BEG2_input[1]),
    .A2(J2MID_ABb_BEG2_input[2]),
    .A3(J2MID_ABb_BEG2_input[3]),
    .S0(ConfigBits[160+0]),
    .S0N(ConfigBits_N[160+0]),
    .S1(ConfigBits[160+1]),
    .S1N(ConfigBits_N[160+1]),
    .X(J2MID_ABb_BEG2)
);

 //switch matrix multiplexer J2MID_ABb_BEG3 MUX-4
assign J2MID_ABb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG3 (
    .A0(J2MID_ABb_BEG3_input[0]),
    .A1(J2MID_ABb_BEG3_input[1]),
    .A2(J2MID_ABb_BEG3_input[2]),
    .A3(J2MID_ABb_BEG3_input[3]),
    .S0(ConfigBits[162+0]),
    .S0N(ConfigBits_N[162+0]),
    .S1(ConfigBits[162+1]),
    .S1N(ConfigBits_N[162+1]),
    .X(J2MID_ABb_BEG3)
);

 //switch matrix multiplexer J2MID_CDb_BEG0 MUX-4
assign J2MID_CDb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG0 (
    .A0(J2MID_CDb_BEG0_input[0]),
    .A1(J2MID_CDb_BEG0_input[1]),
    .A2(J2MID_CDb_BEG0_input[2]),
    .A3(J2MID_CDb_BEG0_input[3]),
    .S0(ConfigBits[164+0]),
    .S0N(ConfigBits_N[164+0]),
    .S1(ConfigBits[164+1]),
    .S1N(ConfigBits_N[164+1]),
    .X(J2MID_CDb_BEG0)
);

 //switch matrix multiplexer J2MID_CDb_BEG1 MUX-4
assign J2MID_CDb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG1 (
    .A0(J2MID_CDb_BEG1_input[0]),
    .A1(J2MID_CDb_BEG1_input[1]),
    .A2(J2MID_CDb_BEG1_input[2]),
    .A3(J2MID_CDb_BEG1_input[3]),
    .S0(ConfigBits[166+0]),
    .S0N(ConfigBits_N[166+0]),
    .S1(ConfigBits[166+1]),
    .S1N(ConfigBits_N[166+1]),
    .X(J2MID_CDb_BEG1)
);

 //switch matrix multiplexer J2MID_CDb_BEG2 MUX-4
assign J2MID_CDb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG2 (
    .A0(J2MID_CDb_BEG2_input[0]),
    .A1(J2MID_CDb_BEG2_input[1]),
    .A2(J2MID_CDb_BEG2_input[2]),
    .A3(J2MID_CDb_BEG2_input[3]),
    .S0(ConfigBits[168+0]),
    .S0N(ConfigBits_N[168+0]),
    .S1(ConfigBits[168+1]),
    .S1N(ConfigBits_N[168+1]),
    .X(J2MID_CDb_BEG2)
);

 //switch matrix multiplexer J2MID_CDb_BEG3 MUX-4
assign J2MID_CDb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG3 (
    .A0(J2MID_CDb_BEG3_input[0]),
    .A1(J2MID_CDb_BEG3_input[1]),
    .A2(J2MID_CDb_BEG3_input[2]),
    .A3(J2MID_CDb_BEG3_input[3]),
    .S0(ConfigBits[170+0]),
    .S0N(ConfigBits_N[170+0]),
    .S1(ConfigBits[170+1]),
    .S1N(ConfigBits_N[170+1]),
    .X(J2MID_CDb_BEG3)
);

 //switch matrix multiplexer J2MID_EFb_BEG0 MUX-4
assign J2MID_EFb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG0 (
    .A0(J2MID_EFb_BEG0_input[0]),
    .A1(J2MID_EFb_BEG0_input[1]),
    .A2(J2MID_EFb_BEG0_input[2]),
    .A3(J2MID_EFb_BEG0_input[3]),
    .S0(ConfigBits[172+0]),
    .S0N(ConfigBits_N[172+0]),
    .S1(ConfigBits[172+1]),
    .S1N(ConfigBits_N[172+1]),
    .X(J2MID_EFb_BEG0)
);

 //switch matrix multiplexer J2MID_EFb_BEG1 MUX-4
assign J2MID_EFb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG1 (
    .A0(J2MID_EFb_BEG1_input[0]),
    .A1(J2MID_EFb_BEG1_input[1]),
    .A2(J2MID_EFb_BEG1_input[2]),
    .A3(J2MID_EFb_BEG1_input[3]),
    .S0(ConfigBits[174+0]),
    .S0N(ConfigBits_N[174+0]),
    .S1(ConfigBits[174+1]),
    .S1N(ConfigBits_N[174+1]),
    .X(J2MID_EFb_BEG1)
);

 //switch matrix multiplexer J2MID_EFb_BEG2 MUX-4
assign J2MID_EFb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG2 (
    .A0(J2MID_EFb_BEG2_input[0]),
    .A1(J2MID_EFb_BEG2_input[1]),
    .A2(J2MID_EFb_BEG2_input[2]),
    .A3(J2MID_EFb_BEG2_input[3]),
    .S0(ConfigBits[176+0]),
    .S0N(ConfigBits_N[176+0]),
    .S1(ConfigBits[176+1]),
    .S1N(ConfigBits_N[176+1]),
    .X(J2MID_EFb_BEG2)
);

 //switch matrix multiplexer J2MID_EFb_BEG3 MUX-4
assign J2MID_EFb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG3 (
    .A0(J2MID_EFb_BEG3_input[0]),
    .A1(J2MID_EFb_BEG3_input[1]),
    .A2(J2MID_EFb_BEG3_input[2]),
    .A3(J2MID_EFb_BEG3_input[3]),
    .S0(ConfigBits[178+0]),
    .S0N(ConfigBits_N[178+0]),
    .S1(ConfigBits[178+1]),
    .S1N(ConfigBits_N[178+1]),
    .X(J2MID_EFb_BEG3)
);

 //switch matrix multiplexer J2MID_GHb_BEG0 MUX-4
assign J2MID_GHb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG0 (
    .A0(J2MID_GHb_BEG0_input[0]),
    .A1(J2MID_GHb_BEG0_input[1]),
    .A2(J2MID_GHb_BEG0_input[2]),
    .A3(J2MID_GHb_BEG0_input[3]),
    .S0(ConfigBits[180+0]),
    .S0N(ConfigBits_N[180+0]),
    .S1(ConfigBits[180+1]),
    .S1N(ConfigBits_N[180+1]),
    .X(J2MID_GHb_BEG0)
);

 //switch matrix multiplexer J2MID_GHb_BEG1 MUX-4
assign J2MID_GHb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG1 (
    .A0(J2MID_GHb_BEG1_input[0]),
    .A1(J2MID_GHb_BEG1_input[1]),
    .A2(J2MID_GHb_BEG1_input[2]),
    .A3(J2MID_GHb_BEG1_input[3]),
    .S0(ConfigBits[182+0]),
    .S0N(ConfigBits_N[182+0]),
    .S1(ConfigBits[182+1]),
    .S1N(ConfigBits_N[182+1]),
    .X(J2MID_GHb_BEG1)
);

 //switch matrix multiplexer J2MID_GHb_BEG2 MUX-4
assign J2MID_GHb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG2 (
    .A0(J2MID_GHb_BEG2_input[0]),
    .A1(J2MID_GHb_BEG2_input[1]),
    .A2(J2MID_GHb_BEG2_input[2]),
    .A3(J2MID_GHb_BEG2_input[3]),
    .S0(ConfigBits[184+0]),
    .S0N(ConfigBits_N[184+0]),
    .S1(ConfigBits[184+1]),
    .S1N(ConfigBits_N[184+1]),
    .X(J2MID_GHb_BEG2)
);

 //switch matrix multiplexer J2MID_GHb_BEG3 MUX-4
assign J2MID_GHb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG3 (
    .A0(J2MID_GHb_BEG3_input[0]),
    .A1(J2MID_GHb_BEG3_input[1]),
    .A2(J2MID_GHb_BEG3_input[2]),
    .A3(J2MID_GHb_BEG3_input[3]),
    .S0(ConfigBits[186+0]),
    .S0N(ConfigBits_N[186+0]),
    .S1(ConfigBits[186+1]),
    .S1N(ConfigBits_N[186+1]),
    .X(J2MID_GHb_BEG3)
);

 //switch matrix multiplexer J2END_AB_BEG0 MUX-4
assign J2END_AB_BEG0_input = {W2END6,SS4END3,E2END6,N2END6};
cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG0 (
    .A0(J2END_AB_BEG0_input[0]),
    .A1(J2END_AB_BEG0_input[1]),
    .A2(J2END_AB_BEG0_input[2]),
    .A3(J2END_AB_BEG0_input[3]),
    .S0(ConfigBits[188+0]),
    .S0N(ConfigBits_N[188+0]),
    .S1(ConfigBits[188+1]),
    .S1N(ConfigBits_N[188+1]),
    .X(J2END_AB_BEG0)
);

 //switch matrix multiplexer J2END_AB_BEG1 MUX-4
assign J2END_AB_BEG1_input = {W2END2,S2END2,E2END2,NN4END0};
cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG1 (
    .A0(J2END_AB_BEG1_input[0]),
    .A1(J2END_AB_BEG1_input[1]),
    .A2(J2END_AB_BEG1_input[2]),
    .A3(J2END_AB_BEG1_input[3]),
    .S0(ConfigBits[190+0]),
    .S0N(ConfigBits_N[190+0]),
    .S1(ConfigBits[190+1]),
    .S1N(ConfigBits_N[190+1]),
    .X(J2END_AB_BEG1)
);

 //switch matrix multiplexer J2END_AB_BEG2 MUX-4
assign J2END_AB_BEG2_input = {W2END4,S2END4,EE4END0,N2END4};
cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG2 (
    .A0(J2END_AB_BEG2_input[0]),
    .A1(J2END_AB_BEG2_input[1]),
    .A2(J2END_AB_BEG2_input[2]),
    .A3(J2END_AB_BEG2_input[3]),
    .S0(ConfigBits[192+0]),
    .S0N(ConfigBits_N[192+0]),
    .S1(ConfigBits[192+1]),
    .S1N(ConfigBits_N[192+1]),
    .X(J2END_AB_BEG2)
);

 //switch matrix multiplexer J2END_AB_BEG3 MUX-4
assign J2END_AB_BEG3_input = {WW4END3,S2END0,E2END0,N2END0};
cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG3 (
    .A0(J2END_AB_BEG3_input[0]),
    .A1(J2END_AB_BEG3_input[1]),
    .A2(J2END_AB_BEG3_input[2]),
    .A3(J2END_AB_BEG3_input[3]),
    .S0(ConfigBits[194+0]),
    .S0N(ConfigBits_N[194+0]),
    .S1(ConfigBits[194+1]),
    .S1N(ConfigBits_N[194+1]),
    .X(J2END_AB_BEG3)
);

 //switch matrix multiplexer J2END_CD_BEG0 MUX-4
assign J2END_CD_BEG0_input = {W2END6,S2END6,E2END6,NN4END3};
cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG0 (
    .A0(J2END_CD_BEG0_input[0]),
    .A1(J2END_CD_BEG0_input[1]),
    .A2(J2END_CD_BEG0_input[2]),
    .A3(J2END_CD_BEG0_input[3]),
    .S0(ConfigBits[196+0]),
    .S0N(ConfigBits_N[196+0]),
    .S1(ConfigBits[196+1]),
    .S1N(ConfigBits_N[196+1]),
    .X(J2END_CD_BEG0)
);

 //switch matrix multiplexer J2END_CD_BEG1 MUX-4
assign J2END_CD_BEG1_input = {WW4END2,S2END2,E2END2,N2END2};
cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG1 (
    .A0(J2END_CD_BEG1_input[0]),
    .A1(J2END_CD_BEG1_input[1]),
    .A2(J2END_CD_BEG1_input[2]),
    .A3(J2END_CD_BEG1_input[3]),
    .S0(ConfigBits[198+0]),
    .S0N(ConfigBits_N[198+0]),
    .S1(ConfigBits[198+1]),
    .S1N(ConfigBits_N[198+1]),
    .X(J2END_CD_BEG1)
);

 //switch matrix multiplexer J2END_CD_BEG2 MUX-4
assign J2END_CD_BEG2_input = {W2END4,SS4END2,E2END4,N2END4};
cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG2 (
    .A0(J2END_CD_BEG2_input[0]),
    .A1(J2END_CD_BEG2_input[1]),
    .A2(J2END_CD_BEG2_input[2]),
    .A3(J2END_CD_BEG2_input[3]),
    .S0(ConfigBits[200+0]),
    .S0N(ConfigBits_N[200+0]),
    .S1(ConfigBits[200+1]),
    .S1N(ConfigBits_N[200+1]),
    .X(J2END_CD_BEG2)
);

 //switch matrix multiplexer J2END_CD_BEG3 MUX-4
assign J2END_CD_BEG3_input = {W2END0,S2END0,EE4END1,N2END0};
cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG3 (
    .A0(J2END_CD_BEG3_input[0]),
    .A1(J2END_CD_BEG3_input[1]),
    .A2(J2END_CD_BEG3_input[2]),
    .A3(J2END_CD_BEG3_input[3]),
    .S0(ConfigBits[202+0]),
    .S0N(ConfigBits_N[202+0]),
    .S1(ConfigBits[202+1]),
    .S1N(ConfigBits_N[202+1]),
    .X(J2END_CD_BEG3)
);

 //switch matrix multiplexer J2END_EF_BEG0 MUX-4
assign J2END_EF_BEG0_input = {W2END7,S2END7,EE4END2,N2END7};
cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG0 (
    .A0(J2END_EF_BEG0_input[0]),
    .A1(J2END_EF_BEG0_input[1]),
    .A2(J2END_EF_BEG0_input[2]),
    .A3(J2END_EF_BEG0_input[3]),
    .S0(ConfigBits[204+0]),
    .S0N(ConfigBits_N[204+0]),
    .S1(ConfigBits[204+1]),
    .S1N(ConfigBits_N[204+1]),
    .X(J2END_EF_BEG0)
);

 //switch matrix multiplexer J2END_EF_BEG1 MUX-4
assign J2END_EF_BEG1_input = {WW4END1,S2END3,E2END3,N2END3};
cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG1 (
    .A0(J2END_EF_BEG1_input[0]),
    .A1(J2END_EF_BEG1_input[1]),
    .A2(J2END_EF_BEG1_input[2]),
    .A3(J2END_EF_BEG1_input[3]),
    .S0(ConfigBits[206+0]),
    .S0N(ConfigBits_N[206+0]),
    .S1(ConfigBits[206+1]),
    .S1N(ConfigBits_N[206+1]),
    .X(J2END_EF_BEG1)
);

 //switch matrix multiplexer J2END_EF_BEG2 MUX-4
assign J2END_EF_BEG2_input = {W2END5,SS4END1,E2END5,N2END5};
cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG2 (
    .A0(J2END_EF_BEG2_input[0]),
    .A1(J2END_EF_BEG2_input[1]),
    .A2(J2END_EF_BEG2_input[2]),
    .A3(J2END_EF_BEG2_input[3]),
    .S0(ConfigBits[208+0]),
    .S0N(ConfigBits_N[208+0]),
    .S1(ConfigBits[208+1]),
    .S1N(ConfigBits_N[208+1]),
    .X(J2END_EF_BEG2)
);

 //switch matrix multiplexer J2END_EF_BEG3 MUX-4
assign J2END_EF_BEG3_input = {W2END1,S2END1,E2END1,NN4END2};
cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG3 (
    .A0(J2END_EF_BEG3_input[0]),
    .A1(J2END_EF_BEG3_input[1]),
    .A2(J2END_EF_BEG3_input[2]),
    .A3(J2END_EF_BEG3_input[3]),
    .S0(ConfigBits[210+0]),
    .S0N(ConfigBits_N[210+0]),
    .S1(ConfigBits[210+1]),
    .S1N(ConfigBits_N[210+1]),
    .X(J2END_EF_BEG3)
);

 //switch matrix multiplexer J2END_GH_BEG0 MUX-4
assign J2END_GH_BEG0_input = {WW4END0,S2END7,E2END7,N2END7};
cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG0 (
    .A0(J2END_GH_BEG0_input[0]),
    .A1(J2END_GH_BEG0_input[1]),
    .A2(J2END_GH_BEG0_input[2]),
    .A3(J2END_GH_BEG0_input[3]),
    .S0(ConfigBits[212+0]),
    .S0N(ConfigBits_N[212+0]),
    .S1(ConfigBits[212+1]),
    .S1N(ConfigBits_N[212+1]),
    .X(J2END_GH_BEG0)
);

 //switch matrix multiplexer J2END_GH_BEG1 MUX-4
assign J2END_GH_BEG1_input = {W2END3,SS4END0,E2END3,N2END3};
cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG1 (
    .A0(J2END_GH_BEG1_input[0]),
    .A1(J2END_GH_BEG1_input[1]),
    .A2(J2END_GH_BEG1_input[2]),
    .A3(J2END_GH_BEG1_input[3]),
    .S0(ConfigBits[214+0]),
    .S0N(ConfigBits_N[214+0]),
    .S1(ConfigBits[214+1]),
    .S1N(ConfigBits_N[214+1]),
    .X(J2END_GH_BEG1)
);

 //switch matrix multiplexer J2END_GH_BEG2 MUX-4
assign J2END_GH_BEG2_input = {W2END5,S2END5,E2END5,NN4END1};
cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG2 (
    .A0(J2END_GH_BEG2_input[0]),
    .A1(J2END_GH_BEG2_input[1]),
    .A2(J2END_GH_BEG2_input[2]),
    .A3(J2END_GH_BEG2_input[3]),
    .S0(ConfigBits[216+0]),
    .S0N(ConfigBits_N[216+0]),
    .S1(ConfigBits[216+1]),
    .S1N(ConfigBits_N[216+1]),
    .X(J2END_GH_BEG2)
);

 //switch matrix multiplexer J2END_GH_BEG3 MUX-4
assign J2END_GH_BEG3_input = {W2END1,S2END1,EE4END3,N2END1};
cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG3 (
    .A0(J2END_GH_BEG3_input[0]),
    .A1(J2END_GH_BEG3_input[1]),
    .A2(J2END_GH_BEG3_input[2]),
    .A3(J2END_GH_BEG3_input[3]),
    .S0(ConfigBits[218+0]),
    .S0N(ConfigBits_N[218+0]),
    .S1(ConfigBits[218+1]),
    .S1N(ConfigBits_N[218+1]),
    .X(J2END_GH_BEG3)
);

 //switch matrix multiplexer JN2BEG0 MUX-16
assign JN2BEG0_input = {resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W6END1,W2END1,S4END1,S4END0,S2END1,E6END1,EE4END0,E2END1,E1END3,N4END1,N2END1};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG0 (
    .A0(JN2BEG0_input[0]),
    .A1(JN2BEG0_input[1]),
    .A2(JN2BEG0_input[2]),
    .A3(JN2BEG0_input[3]),
    .A4(JN2BEG0_input[4]),
    .A5(JN2BEG0_input[5]),
    .A6(JN2BEG0_input[6]),
    .A7(JN2BEG0_input[7]),
    .A8(JN2BEG0_input[8]),
    .A9(JN2BEG0_input[9]),
    .A10(JN2BEG0_input[10]),
    .A11(JN2BEG0_input[11]),
    .A12(JN2BEG0_input[12]),
    .A13(JN2BEG0_input[13]),
    .A14(JN2BEG0_input[14]),
    .A15(JN2BEG0_input[15]),
    .S0(ConfigBits[220+0]),
    .S0N(ConfigBits_N[220+0]),
    .S1(ConfigBits[220+1]),
    .S1N(ConfigBits_N[220+1]),
    .S2(ConfigBits[220+2]),
    .S2N(ConfigBits_N[220+2]),
    .S3(ConfigBits[220+3]),
    .S3N(ConfigBits_N[220+3]),
    .X(JN2BEG0)
);

 //switch matrix multiplexer JN2BEG1 MUX-16
assign JN2BEG1_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,W6END0,W2END2,S4END1,S4END0,S2END2,E6END0,EE4END1,E2END2,E1END0,N4END2,N2END2};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG1 (
    .A0(JN2BEG1_input[0]),
    .A1(JN2BEG1_input[1]),
    .A2(JN2BEG1_input[2]),
    .A3(JN2BEG1_input[3]),
    .A4(JN2BEG1_input[4]),
    .A5(JN2BEG1_input[5]),
    .A6(JN2BEG1_input[6]),
    .A7(JN2BEG1_input[7]),
    .A8(JN2BEG1_input[8]),
    .A9(JN2BEG1_input[9]),
    .A10(JN2BEG1_input[10]),
    .A11(JN2BEG1_input[11]),
    .A12(JN2BEG1_input[12]),
    .A13(JN2BEG1_input[13]),
    .A14(JN2BEG1_input[14]),
    .A15(JN2BEG1_input[15]),
    .S0(ConfigBits[224+0]),
    .S0N(ConfigBits_N[224+0]),
    .S1(ConfigBits[224+1]),
    .S1N(ConfigBits_N[224+1]),
    .S2(ConfigBits[224+2]),
    .S2N(ConfigBits_N[224+2]),
    .S3(ConfigBits[224+3]),
    .S3N(ConfigBits_N[224+3]),
    .X(JN2BEG1)
);

 //switch matrix multiplexer JN2BEG2 MUX-16
assign JN2BEG2_input = {t_resp_ready,resp_status2,resp_status1,resp_status0,req_ready,W6END1,WW4END2,W2END3,S4END1,S4END0,S2END3,E6END1,E2END3,E1END1,N4END3,N2END3};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG2 (
    .A0(JN2BEG2_input[0]),
    .A1(JN2BEG2_input[1]),
    .A2(JN2BEG2_input[2]),
    .A3(JN2BEG2_input[3]),
    .A4(JN2BEG2_input[4]),
    .A5(JN2BEG2_input[5]),
    .A6(JN2BEG2_input[6]),
    .A7(JN2BEG2_input[7]),
    .A8(JN2BEG2_input[8]),
    .A9(JN2BEG2_input[9]),
    .A10(JN2BEG2_input[10]),
    .A11(JN2BEG2_input[11]),
    .A12(JN2BEG2_input[12]),
    .A13(JN2BEG2_input[13]),
    .A14(JN2BEG2_input[14]),
    .A15(JN2BEG2_input[15]),
    .S0(ConfigBits[228+0]),
    .S0N(ConfigBits_N[228+0]),
    .S1(ConfigBits[228+1]),
    .S1N(ConfigBits_N[228+1]),
    .S2(ConfigBits[228+2]),
    .S2N(ConfigBits_N[228+2]),
    .S3(ConfigBits[228+3]),
    .S3N(ConfigBits_N[228+3]),
    .X(JN2BEG2)
);

 //switch matrix multiplexer JN2BEG3 MUX-16
assign JN2BEG3_input = {t_resp_ready,resp_valid,resp_status1,resp_status0,req_ready,W6END0,WW4END3,W2END4,S4END1,S4END0,S2END4,E6END0,E2END4,E1END2,N4END0,N2END4};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG3 (
    .A0(JN2BEG3_input[0]),
    .A1(JN2BEG3_input[1]),
    .A2(JN2BEG3_input[2]),
    .A3(JN2BEG3_input[3]),
    .A4(JN2BEG3_input[4]),
    .A5(JN2BEG3_input[5]),
    .A6(JN2BEG3_input[6]),
    .A7(JN2BEG3_input[7]),
    .A8(JN2BEG3_input[8]),
    .A9(JN2BEG3_input[9]),
    .A10(JN2BEG3_input[10]),
    .A11(JN2BEG3_input[11]),
    .A12(JN2BEG3_input[12]),
    .A13(JN2BEG3_input[13]),
    .A14(JN2BEG3_input[14]),
    .A15(JN2BEG3_input[15]),
    .S0(ConfigBits[232+0]),
    .S0N(ConfigBits_N[232+0]),
    .S1(ConfigBits[232+1]),
    .S1N(ConfigBits_N[232+1]),
    .S2(ConfigBits[232+2]),
    .S2N(ConfigBits_N[232+2]),
    .S3(ConfigBits[232+3]),
    .S3N(ConfigBits_N[232+3]),
    .X(JN2BEG3)
);

 //switch matrix multiplexer JN2BEG4 MUX-16
assign JN2BEG4_input = {t_resp_ready,resp_valid,resp_status2,resp_status0,req_ready,W1END3,W1END1,S4END1,S4END0,S2END5,S1END1,E2END5,E1END1,NN4END3,N2END5,N1END1};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG4 (
    .A0(JN2BEG4_input[0]),
    .A1(JN2BEG4_input[1]),
    .A2(JN2BEG4_input[2]),
    .A3(JN2BEG4_input[3]),
    .A4(JN2BEG4_input[4]),
    .A5(JN2BEG4_input[5]),
    .A6(JN2BEG4_input[6]),
    .A7(JN2BEG4_input[7]),
    .A8(JN2BEG4_input[8]),
    .A9(JN2BEG4_input[9]),
    .A10(JN2BEG4_input[10]),
    .A11(JN2BEG4_input[11]),
    .A12(JN2BEG4_input[12]),
    .A13(JN2BEG4_input[13]),
    .A14(JN2BEG4_input[14]),
    .A15(JN2BEG4_input[15]),
    .S0(ConfigBits[236+0]),
    .S0N(ConfigBits_N[236+0]),
    .S1(ConfigBits[236+1]),
    .S1N(ConfigBits_N[236+1]),
    .S2(ConfigBits[236+2]),
    .S2N(ConfigBits_N[236+2]),
    .S3(ConfigBits[236+3]),
    .S3N(ConfigBits_N[236+3]),
    .X(JN2BEG4)
);

 //switch matrix multiplexer JN2BEG5 MUX-16
assign JN2BEG5_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,req_ready,W1END2,W1END0,S4END1,S4END0,S2END6,S1END2,E2END6,E1END2,NN4END2,N2END6,N1END2};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG5 (
    .A0(JN2BEG5_input[0]),
    .A1(JN2BEG5_input[1]),
    .A2(JN2BEG5_input[2]),
    .A3(JN2BEG5_input[3]),
    .A4(JN2BEG5_input[4]),
    .A5(JN2BEG5_input[5]),
    .A6(JN2BEG5_input[6]),
    .A7(JN2BEG5_input[7]),
    .A8(JN2BEG5_input[8]),
    .A9(JN2BEG5_input[9]),
    .A10(JN2BEG5_input[10]),
    .A11(JN2BEG5_input[11]),
    .A12(JN2BEG5_input[12]),
    .A13(JN2BEG5_input[13]),
    .A14(JN2BEG5_input[14]),
    .A15(JN2BEG5_input[15]),
    .S0(ConfigBits[240+0]),
    .S0N(ConfigBits_N[240+0]),
    .S1(ConfigBits[240+1]),
    .S1N(ConfigBits_N[240+1]),
    .S2(ConfigBits[240+2]),
    .S2N(ConfigBits_N[240+2]),
    .S3(ConfigBits[240+3]),
    .S3N(ConfigBits_N[240+3]),
    .X(JN2BEG5)
);

 //switch matrix multiplexer JN2BEG6 MUX-16
assign JN2BEG6_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END3,W1END1,S4END1,S2END7,S1END3,E2END7,E1END3,NN4END1,N2END7,N1END3};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG6 (
    .A0(JN2BEG6_input[0]),
    .A1(JN2BEG6_input[1]),
    .A2(JN2BEG6_input[2]),
    .A3(JN2BEG6_input[3]),
    .A4(JN2BEG6_input[4]),
    .A5(JN2BEG6_input[5]),
    .A6(JN2BEG6_input[6]),
    .A7(JN2BEG6_input[7]),
    .A8(JN2BEG6_input[8]),
    .A9(JN2BEG6_input[9]),
    .A10(JN2BEG6_input[10]),
    .A11(JN2BEG6_input[11]),
    .A12(JN2BEG6_input[12]),
    .A13(JN2BEG6_input[13]),
    .A14(JN2BEG6_input[14]),
    .A15(JN2BEG6_input[15]),
    .S0(ConfigBits[244+0]),
    .S0N(ConfigBits_N[244+0]),
    .S1(ConfigBits[244+1]),
    .S1N(ConfigBits_N[244+1]),
    .S2(ConfigBits[244+2]),
    .S2N(ConfigBits_N[244+2]),
    .S3(ConfigBits[244+3]),
    .S3N(ConfigBits_N[244+3]),
    .X(JN2BEG6)
);

 //switch matrix multiplexer JN2BEG7 MUX-16
assign JN2BEG7_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END2,W1END0,S4END0,S2END0,S1END0,E2END0,E1END0,NN4END0,N2END0,N1END0};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG7 (
    .A0(JN2BEG7_input[0]),
    .A1(JN2BEG7_input[1]),
    .A2(JN2BEG7_input[2]),
    .A3(JN2BEG7_input[3]),
    .A4(JN2BEG7_input[4]),
    .A5(JN2BEG7_input[5]),
    .A6(JN2BEG7_input[6]),
    .A7(JN2BEG7_input[7]),
    .A8(JN2BEG7_input[8]),
    .A9(JN2BEG7_input[9]),
    .A10(JN2BEG7_input[10]),
    .A11(JN2BEG7_input[11]),
    .A12(JN2BEG7_input[12]),
    .A13(JN2BEG7_input[13]),
    .A14(JN2BEG7_input[14]),
    .A15(JN2BEG7_input[15]),
    .S0(ConfigBits[248+0]),
    .S0N(ConfigBits_N[248+0]),
    .S1(ConfigBits[248+1]),
    .S1N(ConfigBits_N[248+1]),
    .S2(ConfigBits[248+2]),
    .S2N(ConfigBits_N[248+2]),
    .S3(ConfigBits[248+3]),
    .S3N(ConfigBits_N[248+3]),
    .X(JN2BEG7)
);

 //switch matrix multiplexer JE2BEG0 MUX-16
assign JE2BEG0_input = {resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W6END1,W2END1,S4END1,S4END0,S2END1,E6END1,E2END1,NN4END0,N4END1,N2END1,N1END3};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG0 (
    .A0(JE2BEG0_input[0]),
    .A1(JE2BEG0_input[1]),
    .A2(JE2BEG0_input[2]),
    .A3(JE2BEG0_input[3]),
    .A4(JE2BEG0_input[4]),
    .A5(JE2BEG0_input[5]),
    .A6(JE2BEG0_input[6]),
    .A7(JE2BEG0_input[7]),
    .A8(JE2BEG0_input[8]),
    .A9(JE2BEG0_input[9]),
    .A10(JE2BEG0_input[10]),
    .A11(JE2BEG0_input[11]),
    .A12(JE2BEG0_input[12]),
    .A13(JE2BEG0_input[13]),
    .A14(JE2BEG0_input[14]),
    .A15(JE2BEG0_input[15]),
    .S0(ConfigBits[252+0]),
    .S0N(ConfigBits_N[252+0]),
    .S1(ConfigBits[252+1]),
    .S1N(ConfigBits_N[252+1]),
    .S2(ConfigBits[252+2]),
    .S2N(ConfigBits_N[252+2]),
    .S3(ConfigBits[252+3]),
    .S3N(ConfigBits_N[252+3]),
    .X(JE2BEG0)
);

 //switch matrix multiplexer JE2BEG1 MUX-16
assign JE2BEG1_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,W6END0,W2END2,S4END1,S4END0,S2END2,E6END0,E2END2,NN4END1,N4END2,N2END2,N1END0};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG1 (
    .A0(JE2BEG1_input[0]),
    .A1(JE2BEG1_input[1]),
    .A2(JE2BEG1_input[2]),
    .A3(JE2BEG1_input[3]),
    .A4(JE2BEG1_input[4]),
    .A5(JE2BEG1_input[5]),
    .A6(JE2BEG1_input[6]),
    .A7(JE2BEG1_input[7]),
    .A8(JE2BEG1_input[8]),
    .A9(JE2BEG1_input[9]),
    .A10(JE2BEG1_input[10]),
    .A11(JE2BEG1_input[11]),
    .A12(JE2BEG1_input[12]),
    .A13(JE2BEG1_input[13]),
    .A14(JE2BEG1_input[14]),
    .A15(JE2BEG1_input[15]),
    .S0(ConfigBits[256+0]),
    .S0N(ConfigBits_N[256+0]),
    .S1(ConfigBits[256+1]),
    .S1N(ConfigBits_N[256+1]),
    .S2(ConfigBits[256+2]),
    .S2N(ConfigBits_N[256+2]),
    .S3(ConfigBits[256+3]),
    .S3N(ConfigBits_N[256+3]),
    .X(JE2BEG1)
);

 //switch matrix multiplexer JE2BEG2 MUX-16
assign JE2BEG2_input = {t_resp_ready,resp_status2,resp_status1,resp_status0,req_ready,W6END1,W2END3,SS4END2,S4END1,S4END0,S2END3,E6END1,E2END3,N4END3,N2END3,N1END1};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG2 (
    .A0(JE2BEG2_input[0]),
    .A1(JE2BEG2_input[1]),
    .A2(JE2BEG2_input[2]),
    .A3(JE2BEG2_input[3]),
    .A4(JE2BEG2_input[4]),
    .A5(JE2BEG2_input[5]),
    .A6(JE2BEG2_input[6]),
    .A7(JE2BEG2_input[7]),
    .A8(JE2BEG2_input[8]),
    .A9(JE2BEG2_input[9]),
    .A10(JE2BEG2_input[10]),
    .A11(JE2BEG2_input[11]),
    .A12(JE2BEG2_input[12]),
    .A13(JE2BEG2_input[13]),
    .A14(JE2BEG2_input[14]),
    .A15(JE2BEG2_input[15]),
    .S0(ConfigBits[260+0]),
    .S0N(ConfigBits_N[260+0]),
    .S1(ConfigBits[260+1]),
    .S1N(ConfigBits_N[260+1]),
    .S2(ConfigBits[260+2]),
    .S2N(ConfigBits_N[260+2]),
    .S3(ConfigBits[260+3]),
    .S3N(ConfigBits_N[260+3]),
    .X(JE2BEG2)
);

 //switch matrix multiplexer JE2BEG3 MUX-16
assign JE2BEG3_input = {t_resp_ready,resp_valid,resp_status1,resp_status0,req_ready,W6END0,W2END4,SS4END3,S4END1,S4END0,S2END4,E6END0,E2END4,N4END0,N2END4,N1END2};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG3 (
    .A0(JE2BEG3_input[0]),
    .A1(JE2BEG3_input[1]),
    .A2(JE2BEG3_input[2]),
    .A3(JE2BEG3_input[3]),
    .A4(JE2BEG3_input[4]),
    .A5(JE2BEG3_input[5]),
    .A6(JE2BEG3_input[6]),
    .A7(JE2BEG3_input[7]),
    .A8(JE2BEG3_input[8]),
    .A9(JE2BEG3_input[9]),
    .A10(JE2BEG3_input[10]),
    .A11(JE2BEG3_input[11]),
    .A12(JE2BEG3_input[12]),
    .A13(JE2BEG3_input[13]),
    .A14(JE2BEG3_input[14]),
    .A15(JE2BEG3_input[15]),
    .S0(ConfigBits[264+0]),
    .S0N(ConfigBits_N[264+0]),
    .S1(ConfigBits[264+1]),
    .S1N(ConfigBits_N[264+1]),
    .S2(ConfigBits[264+2]),
    .S2N(ConfigBits_N[264+2]),
    .S3(ConfigBits[264+3]),
    .S3N(ConfigBits_N[264+3]),
    .X(JE2BEG3)
);

 //switch matrix multiplexer JE2BEG4 MUX-16
assign JE2BEG4_input = {t_resp_ready,resp_valid,resp_status2,resp_status0,req_ready,W1END1,S4END1,S4END0,S2END5,S1END3,S1END1,EE4END3,E2END5,E1END1,N2END5,N1END1};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG4 (
    .A0(JE2BEG4_input[0]),
    .A1(JE2BEG4_input[1]),
    .A2(JE2BEG4_input[2]),
    .A3(JE2BEG4_input[3]),
    .A4(JE2BEG4_input[4]),
    .A5(JE2BEG4_input[5]),
    .A6(JE2BEG4_input[6]),
    .A7(JE2BEG4_input[7]),
    .A8(JE2BEG4_input[8]),
    .A9(JE2BEG4_input[9]),
    .A10(JE2BEG4_input[10]),
    .A11(JE2BEG4_input[11]),
    .A12(JE2BEG4_input[12]),
    .A13(JE2BEG4_input[13]),
    .A14(JE2BEG4_input[14]),
    .A15(JE2BEG4_input[15]),
    .S0(ConfigBits[268+0]),
    .S0N(ConfigBits_N[268+0]),
    .S1(ConfigBits[268+1]),
    .S1N(ConfigBits_N[268+1]),
    .S2(ConfigBits[268+2]),
    .S2N(ConfigBits_N[268+2]),
    .S3(ConfigBits[268+3]),
    .S3N(ConfigBits_N[268+3]),
    .X(JE2BEG4)
);

 //switch matrix multiplexer JE2BEG5 MUX-16
assign JE2BEG5_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,req_ready,W1END2,S4END1,S4END0,S2END6,S1END2,S1END0,EE4END2,E2END6,E1END2,N2END6,N1END2};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG5 (
    .A0(JE2BEG5_input[0]),
    .A1(JE2BEG5_input[1]),
    .A2(JE2BEG5_input[2]),
    .A3(JE2BEG5_input[3]),
    .A4(JE2BEG5_input[4]),
    .A5(JE2BEG5_input[5]),
    .A6(JE2BEG5_input[6]),
    .A7(JE2BEG5_input[7]),
    .A8(JE2BEG5_input[8]),
    .A9(JE2BEG5_input[9]),
    .A10(JE2BEG5_input[10]),
    .A11(JE2BEG5_input[11]),
    .A12(JE2BEG5_input[12]),
    .A13(JE2BEG5_input[13]),
    .A14(JE2BEG5_input[14]),
    .A15(JE2BEG5_input[15]),
    .S0(ConfigBits[272+0]),
    .S0N(ConfigBits_N[272+0]),
    .S1(ConfigBits[272+1]),
    .S1N(ConfigBits_N[272+1]),
    .S2(ConfigBits[272+2]),
    .S2N(ConfigBits_N[272+2]),
    .S3(ConfigBits[272+3]),
    .S3N(ConfigBits_N[272+3]),
    .X(JE2BEG5)
);

 //switch matrix multiplexer JE2BEG6 MUX-16
assign JE2BEG6_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END3,S4END1,S2END7,S1END3,S1END1,EE4END1,E2END7,E1END3,N2END7,N1END3};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG6 (
    .A0(JE2BEG6_input[0]),
    .A1(JE2BEG6_input[1]),
    .A2(JE2BEG6_input[2]),
    .A3(JE2BEG6_input[3]),
    .A4(JE2BEG6_input[4]),
    .A5(JE2BEG6_input[5]),
    .A6(JE2BEG6_input[6]),
    .A7(JE2BEG6_input[7]),
    .A8(JE2BEG6_input[8]),
    .A9(JE2BEG6_input[9]),
    .A10(JE2BEG6_input[10]),
    .A11(JE2BEG6_input[11]),
    .A12(JE2BEG6_input[12]),
    .A13(JE2BEG6_input[13]),
    .A14(JE2BEG6_input[14]),
    .A15(JE2BEG6_input[15]),
    .S0(ConfigBits[276+0]),
    .S0N(ConfigBits_N[276+0]),
    .S1(ConfigBits[276+1]),
    .S1N(ConfigBits_N[276+1]),
    .S2(ConfigBits[276+2]),
    .S2N(ConfigBits_N[276+2]),
    .S3(ConfigBits[276+3]),
    .S3N(ConfigBits_N[276+3]),
    .X(JE2BEG6)
);

 //switch matrix multiplexer JE2BEG7 MUX-16
assign JE2BEG7_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END0,S4END0,S2END0,S1END2,S1END0,EE4END0,E2END0,E1END0,N2END0,N1END0};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG7 (
    .A0(JE2BEG7_input[0]),
    .A1(JE2BEG7_input[1]),
    .A2(JE2BEG7_input[2]),
    .A3(JE2BEG7_input[3]),
    .A4(JE2BEG7_input[4]),
    .A5(JE2BEG7_input[5]),
    .A6(JE2BEG7_input[6]),
    .A7(JE2BEG7_input[7]),
    .A8(JE2BEG7_input[8]),
    .A9(JE2BEG7_input[9]),
    .A10(JE2BEG7_input[10]),
    .A11(JE2BEG7_input[11]),
    .A12(JE2BEG7_input[12]),
    .A13(JE2BEG7_input[13]),
    .A14(JE2BEG7_input[14]),
    .A15(JE2BEG7_input[15]),
    .S0(ConfigBits[280+0]),
    .S0N(ConfigBits_N[280+0]),
    .S1(ConfigBits[280+1]),
    .S1N(ConfigBits_N[280+1]),
    .S2(ConfigBits[280+2]),
    .S2N(ConfigBits_N[280+2]),
    .S3(ConfigBits[280+3]),
    .S3N(ConfigBits_N[280+3]),
    .X(JE2BEG7)
);

 //switch matrix multiplexer JS2BEG0 MUX-15
assign JS2BEG0_input = {resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W6END1,WW4END0,W2END1,S4END1,S4END0,S2END1,E6END1,E2END1,E1END3,N2END1};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG0 (
    .A0(JS2BEG0_input[0]),
    .A1(JS2BEG0_input[1]),
    .A2(JS2BEG0_input[2]),
    .A3(JS2BEG0_input[3]),
    .A4(JS2BEG0_input[4]),
    .A5(JS2BEG0_input[5]),
    .A6(JS2BEG0_input[6]),
    .A7(JS2BEG0_input[7]),
    .A8(JS2BEG0_input[8]),
    .A9(JS2BEG0_input[9]),
    .A10(JS2BEG0_input[10]),
    .A11(JS2BEG0_input[11]),
    .A12(JS2BEG0_input[12]),
    .A13(JS2BEG0_input[13]),
    .A14(JS2BEG0_input[14]),
    .S0(ConfigBits[284+0]),
    .S0N(ConfigBits_N[284+0]),
    .S1(ConfigBits[284+1]),
    .S1N(ConfigBits_N[284+1]),
    .S2(ConfigBits[284+2]),
    .S2N(ConfigBits_N[284+2]),
    .X(JS2BEG0)
);

 //switch matrix multiplexer JS2BEG1 MUX-16
assign JS2BEG1_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,W6END0,WW4END1,W2END2,S4END2,S4END1,S4END0,S2END2,E6END0,E2END2,E1END0,N2END2};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG1 (
    .A0(JS2BEG1_input[0]),
    .A1(JS2BEG1_input[1]),
    .A2(JS2BEG1_input[2]),
    .A3(JS2BEG1_input[3]),
    .A4(JS2BEG1_input[4]),
    .A5(JS2BEG1_input[5]),
    .A6(JS2BEG1_input[6]),
    .A7(JS2BEG1_input[7]),
    .A8(JS2BEG1_input[8]),
    .A9(JS2BEG1_input[9]),
    .A10(JS2BEG1_input[10]),
    .A11(JS2BEG1_input[11]),
    .A12(JS2BEG1_input[12]),
    .A13(JS2BEG1_input[13]),
    .A14(JS2BEG1_input[14]),
    .A15(JS2BEG1_input[15]),
    .S0(ConfigBits[287+0]),
    .S0N(ConfigBits_N[287+0]),
    .S1(ConfigBits[287+1]),
    .S1N(ConfigBits_N[287+1]),
    .S2(ConfigBits[287+2]),
    .S2N(ConfigBits_N[287+2]),
    .S3(ConfigBits[287+3]),
    .S3N(ConfigBits_N[287+3]),
    .X(JS2BEG1)
);

 //switch matrix multiplexer JS2BEG2 MUX-16
assign JS2BEG2_input = {t_resp_ready,resp_status2,resp_status1,resp_status0,req_ready,W6END1,W2END3,S4END3,S4END1,S4END0,S2END3,E6END1,EE4END2,E2END3,E1END1,N2END3};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG2 (
    .A0(JS2BEG2_input[0]),
    .A1(JS2BEG2_input[1]),
    .A2(JS2BEG2_input[2]),
    .A3(JS2BEG2_input[3]),
    .A4(JS2BEG2_input[4]),
    .A5(JS2BEG2_input[5]),
    .A6(JS2BEG2_input[6]),
    .A7(JS2BEG2_input[7]),
    .A8(JS2BEG2_input[8]),
    .A9(JS2BEG2_input[9]),
    .A10(JS2BEG2_input[10]),
    .A11(JS2BEG2_input[11]),
    .A12(JS2BEG2_input[12]),
    .A13(JS2BEG2_input[13]),
    .A14(JS2BEG2_input[14]),
    .A15(JS2BEG2_input[15]),
    .S0(ConfigBits[291+0]),
    .S0N(ConfigBits_N[291+0]),
    .S1(ConfigBits[291+1]),
    .S1N(ConfigBits_N[291+1]),
    .S2(ConfigBits[291+2]),
    .S2N(ConfigBits_N[291+2]),
    .S3(ConfigBits[291+3]),
    .S3N(ConfigBits_N[291+3]),
    .X(JS2BEG2)
);

 //switch matrix multiplexer JS2BEG3 MUX-15
assign JS2BEG3_input = {t_resp_ready,resp_valid,resp_status1,resp_status0,req_ready,W6END0,W2END4,S4END1,S4END0,S2END4,E6END0,EE4END3,E2END4,E1END2,N2END4};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG3 (
    .A0(JS2BEG3_input[0]),
    .A1(JS2BEG3_input[1]),
    .A2(JS2BEG3_input[2]),
    .A3(JS2BEG3_input[3]),
    .A4(JS2BEG3_input[4]),
    .A5(JS2BEG3_input[5]),
    .A6(JS2BEG3_input[6]),
    .A7(JS2BEG3_input[7]),
    .A8(JS2BEG3_input[8]),
    .A9(JS2BEG3_input[9]),
    .A10(JS2BEG3_input[10]),
    .A11(JS2BEG3_input[11]),
    .A12(JS2BEG3_input[12]),
    .A13(JS2BEG3_input[13]),
    .A14(JS2BEG3_input[14]),
    .S0(ConfigBits[295+0]),
    .S0N(ConfigBits_N[295+0]),
    .S1(ConfigBits[295+1]),
    .S1N(ConfigBits_N[295+1]),
    .S2(ConfigBits[295+2]),
    .S2N(ConfigBits_N[295+2]),
    .X(JS2BEG3)
);

 //switch matrix multiplexer JS2BEG4 MUX-16
assign JS2BEG4_input = {t_resp_ready,resp_valid,resp_status2,resp_status0,req_ready,W1END3,W1END1,SS4END3,S4END1,S4END0,S2END5,S1END1,E2END5,E1END1,N2END5,N1END1};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG4 (
    .A0(JS2BEG4_input[0]),
    .A1(JS2BEG4_input[1]),
    .A2(JS2BEG4_input[2]),
    .A3(JS2BEG4_input[3]),
    .A4(JS2BEG4_input[4]),
    .A5(JS2BEG4_input[5]),
    .A6(JS2BEG4_input[6]),
    .A7(JS2BEG4_input[7]),
    .A8(JS2BEG4_input[8]),
    .A9(JS2BEG4_input[9]),
    .A10(JS2BEG4_input[10]),
    .A11(JS2BEG4_input[11]),
    .A12(JS2BEG4_input[12]),
    .A13(JS2BEG4_input[13]),
    .A14(JS2BEG4_input[14]),
    .A15(JS2BEG4_input[15]),
    .S0(ConfigBits[298+0]),
    .S0N(ConfigBits_N[298+0]),
    .S1(ConfigBits[298+1]),
    .S1N(ConfigBits_N[298+1]),
    .S2(ConfigBits[298+2]),
    .S2N(ConfigBits_N[298+2]),
    .S3(ConfigBits[298+3]),
    .S3N(ConfigBits_N[298+3]),
    .X(JS2BEG4)
);

 //switch matrix multiplexer JS2BEG5 MUX-16
assign JS2BEG5_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,req_ready,W1END2,W1END0,SS4END2,S4END1,S4END0,S2END6,S1END2,E2END6,E1END2,N2END6,N1END2};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG5 (
    .A0(JS2BEG5_input[0]),
    .A1(JS2BEG5_input[1]),
    .A2(JS2BEG5_input[2]),
    .A3(JS2BEG5_input[3]),
    .A4(JS2BEG5_input[4]),
    .A5(JS2BEG5_input[5]),
    .A6(JS2BEG5_input[6]),
    .A7(JS2BEG5_input[7]),
    .A8(JS2BEG5_input[8]),
    .A9(JS2BEG5_input[9]),
    .A10(JS2BEG5_input[10]),
    .A11(JS2BEG5_input[11]),
    .A12(JS2BEG5_input[12]),
    .A13(JS2BEG5_input[13]),
    .A14(JS2BEG5_input[14]),
    .A15(JS2BEG5_input[15]),
    .S0(ConfigBits[302+0]),
    .S0N(ConfigBits_N[302+0]),
    .S1(ConfigBits[302+1]),
    .S1N(ConfigBits_N[302+1]),
    .S2(ConfigBits[302+2]),
    .S2N(ConfigBits_N[302+2]),
    .S3(ConfigBits[302+3]),
    .S3N(ConfigBits_N[302+3]),
    .X(JS2BEG5)
);

 //switch matrix multiplexer JS2BEG6 MUX-16
assign JS2BEG6_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END3,W1END1,SS4END1,S4END1,S2END7,S1END3,E2END7,E1END3,N2END7,N1END3};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG6 (
    .A0(JS2BEG6_input[0]),
    .A1(JS2BEG6_input[1]),
    .A2(JS2BEG6_input[2]),
    .A3(JS2BEG6_input[3]),
    .A4(JS2BEG6_input[4]),
    .A5(JS2BEG6_input[5]),
    .A6(JS2BEG6_input[6]),
    .A7(JS2BEG6_input[7]),
    .A8(JS2BEG6_input[8]),
    .A9(JS2BEG6_input[9]),
    .A10(JS2BEG6_input[10]),
    .A11(JS2BEG6_input[11]),
    .A12(JS2BEG6_input[12]),
    .A13(JS2BEG6_input[13]),
    .A14(JS2BEG6_input[14]),
    .A15(JS2BEG6_input[15]),
    .S0(ConfigBits[306+0]),
    .S0N(ConfigBits_N[306+0]),
    .S1(ConfigBits[306+1]),
    .S1N(ConfigBits_N[306+1]),
    .S2(ConfigBits[306+2]),
    .S2N(ConfigBits_N[306+2]),
    .S3(ConfigBits[306+3]),
    .S3N(ConfigBits_N[306+3]),
    .X(JS2BEG6)
);

 //switch matrix multiplexer JS2BEG7 MUX-16
assign JS2BEG7_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W1END2,W1END0,SS4END0,S4END0,S2END0,S1END0,E2END0,E1END0,N2END0,N1END0};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG7 (
    .A0(JS2BEG7_input[0]),
    .A1(JS2BEG7_input[1]),
    .A2(JS2BEG7_input[2]),
    .A3(JS2BEG7_input[3]),
    .A4(JS2BEG7_input[4]),
    .A5(JS2BEG7_input[5]),
    .A6(JS2BEG7_input[6]),
    .A7(JS2BEG7_input[7]),
    .A8(JS2BEG7_input[8]),
    .A9(JS2BEG7_input[9]),
    .A10(JS2BEG7_input[10]),
    .A11(JS2BEG7_input[11]),
    .A12(JS2BEG7_input[12]),
    .A13(JS2BEG7_input[13]),
    .A14(JS2BEG7_input[14]),
    .A15(JS2BEG7_input[15]),
    .S0(ConfigBits[310+0]),
    .S0N(ConfigBits_N[310+0]),
    .S1(ConfigBits[310+1]),
    .S1N(ConfigBits_N[310+1]),
    .S2(ConfigBits[310+2]),
    .S2N(ConfigBits_N[310+2]),
    .S3(ConfigBits[310+3]),
    .S3N(ConfigBits_N[310+3]),
    .X(JS2BEG7)
);

 //switch matrix multiplexer JW2BEG0 MUX-15
assign JW2BEG0_input = {resp_valid,resp_status2,resp_status1,resp_status0,req_ready,W6END1,W2END1,SS4END0,S4END1,S4END0,S2END1,E6END1,E2END1,N2END1,N1END3};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG0 (
    .A0(JW2BEG0_input[0]),
    .A1(JW2BEG0_input[1]),
    .A2(JW2BEG0_input[2]),
    .A3(JW2BEG0_input[3]),
    .A4(JW2BEG0_input[4]),
    .A5(JW2BEG0_input[5]),
    .A6(JW2BEG0_input[6]),
    .A7(JW2BEG0_input[7]),
    .A8(JW2BEG0_input[8]),
    .A9(JW2BEG0_input[9]),
    .A10(JW2BEG0_input[10]),
    .A11(JW2BEG0_input[11]),
    .A12(JW2BEG0_input[12]),
    .A13(JW2BEG0_input[13]),
    .A14(JW2BEG0_input[14]),
    .S0(ConfigBits[314+0]),
    .S0N(ConfigBits_N[314+0]),
    .S1(ConfigBits[314+1]),
    .S1N(ConfigBits_N[314+1]),
    .S2(ConfigBits[314+2]),
    .S2N(ConfigBits_N[314+2]),
    .X(JW2BEG0)
);

 //switch matrix multiplexer JW2BEG1 MUX-16
assign JW2BEG1_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,W6END0,W2END2,SS4END1,S4END2,S4END1,S4END0,S2END2,E6END0,E2END2,N2END2,N1END0};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG1 (
    .A0(JW2BEG1_input[0]),
    .A1(JW2BEG1_input[1]),
    .A2(JW2BEG1_input[2]),
    .A3(JW2BEG1_input[3]),
    .A4(JW2BEG1_input[4]),
    .A5(JW2BEG1_input[5]),
    .A6(JW2BEG1_input[6]),
    .A7(JW2BEG1_input[7]),
    .A8(JW2BEG1_input[8]),
    .A9(JW2BEG1_input[9]),
    .A10(JW2BEG1_input[10]),
    .A11(JW2BEG1_input[11]),
    .A12(JW2BEG1_input[12]),
    .A13(JW2BEG1_input[13]),
    .A14(JW2BEG1_input[14]),
    .A15(JW2BEG1_input[15]),
    .S0(ConfigBits[317+0]),
    .S0N(ConfigBits_N[317+0]),
    .S1(ConfigBits[317+1]),
    .S1N(ConfigBits_N[317+1]),
    .S2(ConfigBits[317+2]),
    .S2N(ConfigBits_N[317+2]),
    .S3(ConfigBits[317+3]),
    .S3N(ConfigBits_N[317+3]),
    .X(JW2BEG1)
);

 //switch matrix multiplexer JW2BEG2 MUX-16
assign JW2BEG2_input = {t_resp_ready,resp_status2,resp_status1,resp_status0,req_ready,W6END1,W2END3,S4END3,S4END1,S4END0,S2END3,E6END1,E2END3,NN4END2,N2END3,N1END1};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG2 (
    .A0(JW2BEG2_input[0]),
    .A1(JW2BEG2_input[1]),
    .A2(JW2BEG2_input[2]),
    .A3(JW2BEG2_input[3]),
    .A4(JW2BEG2_input[4]),
    .A5(JW2BEG2_input[5]),
    .A6(JW2BEG2_input[6]),
    .A7(JW2BEG2_input[7]),
    .A8(JW2BEG2_input[8]),
    .A9(JW2BEG2_input[9]),
    .A10(JW2BEG2_input[10]),
    .A11(JW2BEG2_input[11]),
    .A12(JW2BEG2_input[12]),
    .A13(JW2BEG2_input[13]),
    .A14(JW2BEG2_input[14]),
    .A15(JW2BEG2_input[15]),
    .S0(ConfigBits[321+0]),
    .S0N(ConfigBits_N[321+0]),
    .S1(ConfigBits[321+1]),
    .S1N(ConfigBits_N[321+1]),
    .S2(ConfigBits[321+2]),
    .S2N(ConfigBits_N[321+2]),
    .S3(ConfigBits[321+3]),
    .S3N(ConfigBits_N[321+3]),
    .X(JW2BEG2)
);

 //switch matrix multiplexer JW2BEG3 MUX-15
assign JW2BEG3_input = {t_resp_ready,resp_valid,resp_status1,resp_status0,req_ready,W6END0,W2END4,S4END1,S4END0,S2END4,E6END0,E2END4,NN4END3,N2END4,N1END2};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG3 (
    .A0(JW2BEG3_input[0]),
    .A1(JW2BEG3_input[1]),
    .A2(JW2BEG3_input[2]),
    .A3(JW2BEG3_input[3]),
    .A4(JW2BEG3_input[4]),
    .A5(JW2BEG3_input[5]),
    .A6(JW2BEG3_input[6]),
    .A7(JW2BEG3_input[7]),
    .A8(JW2BEG3_input[8]),
    .A9(JW2BEG3_input[9]),
    .A10(JW2BEG3_input[10]),
    .A11(JW2BEG3_input[11]),
    .A12(JW2BEG3_input[12]),
    .A13(JW2BEG3_input[13]),
    .A14(JW2BEG3_input[14]),
    .S0(ConfigBits[325+0]),
    .S0N(ConfigBits_N[325+0]),
    .S1(ConfigBits[325+1]),
    .S1N(ConfigBits_N[325+1]),
    .S2(ConfigBits[325+2]),
    .S2N(ConfigBits_N[325+2]),
    .X(JW2BEG3)
);

 //switch matrix multiplexer JW2BEG4 MUX-16
assign JW2BEG4_input = {t_resp_ready,resp_valid,resp_status2,resp_status0,req_ready,WW4END3,W1END1,S4END1,S4END0,S2END5,S1END3,S1END1,E2END5,E1END1,N2END5,N1END1};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG4 (
    .A0(JW2BEG4_input[0]),
    .A1(JW2BEG4_input[1]),
    .A2(JW2BEG4_input[2]),
    .A3(JW2BEG4_input[3]),
    .A4(JW2BEG4_input[4]),
    .A5(JW2BEG4_input[5]),
    .A6(JW2BEG4_input[6]),
    .A7(JW2BEG4_input[7]),
    .A8(JW2BEG4_input[8]),
    .A9(JW2BEG4_input[9]),
    .A10(JW2BEG4_input[10]),
    .A11(JW2BEG4_input[11]),
    .A12(JW2BEG4_input[12]),
    .A13(JW2BEG4_input[13]),
    .A14(JW2BEG4_input[14]),
    .A15(JW2BEG4_input[15]),
    .S0(ConfigBits[328+0]),
    .S0N(ConfigBits_N[328+0]),
    .S1(ConfigBits[328+1]),
    .S1N(ConfigBits_N[328+1]),
    .S2(ConfigBits[328+2]),
    .S2N(ConfigBits_N[328+2]),
    .S3(ConfigBits[328+3]),
    .S3N(ConfigBits_N[328+3]),
    .X(JW2BEG4)
);

 //switch matrix multiplexer JW2BEG5 MUX-16
assign JW2BEG5_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,req_ready,WW4END2,W1END2,S4END1,S4END0,S2END6,S1END2,S1END0,E2END6,E1END2,N2END6,N1END2};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG5 (
    .A0(JW2BEG5_input[0]),
    .A1(JW2BEG5_input[1]),
    .A2(JW2BEG5_input[2]),
    .A3(JW2BEG5_input[3]),
    .A4(JW2BEG5_input[4]),
    .A5(JW2BEG5_input[5]),
    .A6(JW2BEG5_input[6]),
    .A7(JW2BEG5_input[7]),
    .A8(JW2BEG5_input[8]),
    .A9(JW2BEG5_input[9]),
    .A10(JW2BEG5_input[10]),
    .A11(JW2BEG5_input[11]),
    .A12(JW2BEG5_input[12]),
    .A13(JW2BEG5_input[13]),
    .A14(JW2BEG5_input[14]),
    .A15(JW2BEG5_input[15]),
    .S0(ConfigBits[332+0]),
    .S0N(ConfigBits_N[332+0]),
    .S1(ConfigBits[332+1]),
    .S1N(ConfigBits_N[332+1]),
    .S2(ConfigBits[332+2]),
    .S2N(ConfigBits_N[332+2]),
    .S3(ConfigBits[332+3]),
    .S3N(ConfigBits_N[332+3]),
    .X(JW2BEG5)
);

 //switch matrix multiplexer JW2BEG6 MUX-16
assign JW2BEG6_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,WW4END1,W1END3,S4END1,S2END7,S1END3,S1END1,E2END7,E1END3,N2END7,N1END3};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG6 (
    .A0(JW2BEG6_input[0]),
    .A1(JW2BEG6_input[1]),
    .A2(JW2BEG6_input[2]),
    .A3(JW2BEG6_input[3]),
    .A4(JW2BEG6_input[4]),
    .A5(JW2BEG6_input[5]),
    .A6(JW2BEG6_input[6]),
    .A7(JW2BEG6_input[7]),
    .A8(JW2BEG6_input[8]),
    .A9(JW2BEG6_input[9]),
    .A10(JW2BEG6_input[10]),
    .A11(JW2BEG6_input[11]),
    .A12(JW2BEG6_input[12]),
    .A13(JW2BEG6_input[13]),
    .A14(JW2BEG6_input[14]),
    .A15(JW2BEG6_input[15]),
    .S0(ConfigBits[336+0]),
    .S0N(ConfigBits_N[336+0]),
    .S1(ConfigBits[336+1]),
    .S1N(ConfigBits_N[336+1]),
    .S2(ConfigBits[336+2]),
    .S2N(ConfigBits_N[336+2]),
    .S3(ConfigBits[336+3]),
    .S3N(ConfigBits_N[336+3]),
    .X(JW2BEG6)
);

 //switch matrix multiplexer JW2BEG7 MUX-16
assign JW2BEG7_input = {t_resp_ready,resp_valid,resp_status2,resp_status1,resp_status0,req_ready,WW4END0,W1END0,S4END0,S2END0,S1END2,S1END0,E2END0,E1END0,N2END0,N1END0};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG7 (
    .A0(JW2BEG7_input[0]),
    .A1(JW2BEG7_input[1]),
    .A2(JW2BEG7_input[2]),
    .A3(JW2BEG7_input[3]),
    .A4(JW2BEG7_input[4]),
    .A5(JW2BEG7_input[5]),
    .A6(JW2BEG7_input[6]),
    .A7(JW2BEG7_input[7]),
    .A8(JW2BEG7_input[8]),
    .A9(JW2BEG7_input[9]),
    .A10(JW2BEG7_input[10]),
    .A11(JW2BEG7_input[11]),
    .A12(JW2BEG7_input[12]),
    .A13(JW2BEG7_input[13]),
    .A14(JW2BEG7_input[14]),
    .A15(JW2BEG7_input[15]),
    .S0(ConfigBits[340+0]),
    .S0N(ConfigBits_N[340+0]),
    .S1(ConfigBits[340+1]),
    .S1N(ConfigBits_N[340+1]),
    .S2(ConfigBits[340+2]),
    .S2N(ConfigBits_N[340+2]),
    .S3(ConfigBits[340+3]),
    .S3N(ConfigBits_N[340+3]),
    .X(JW2BEG7)
);

 //switch matrix multiplexer J_l_AB_BEG0 MUX-4
assign J_l_AB_BEG0_input = {JN2END1,WW4END0,S4END3,NN4END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG0 (
    .A0(J_l_AB_BEG0_input[0]),
    .A1(J_l_AB_BEG0_input[1]),
    .A2(J_l_AB_BEG0_input[2]),
    .A3(J_l_AB_BEG0_input[3]),
    .S0(ConfigBits[344+0]),
    .S0N(ConfigBits_N[344+0]),
    .S1(ConfigBits[344+1]),
    .S1N(ConfigBits_N[344+1]),
    .X(J_l_AB_BEG0)
);

 //switch matrix multiplexer J_l_AB_BEG1 MUX-4
assign J_l_AB_BEG1_input = {JE2END1,W2END7,S4END2,EE4END2};
cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG1 (
    .A0(J_l_AB_BEG1_input[0]),
    .A1(J_l_AB_BEG1_input[1]),
    .A2(J_l_AB_BEG1_input[2]),
    .A3(J_l_AB_BEG1_input[3]),
    .S0(ConfigBits[346+0]),
    .S0N(ConfigBits_N[346+0]),
    .S1(ConfigBits[346+1]),
    .S1N(ConfigBits_N[346+1]),
    .X(J_l_AB_BEG1)
);

 //switch matrix multiplexer J_l_AB_BEG2 MUX-4
assign J_l_AB_BEG2_input = {JS2END1,W6END1,E6END1,N4END1};
cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG2 (
    .A0(J_l_AB_BEG2_input[0]),
    .A1(J_l_AB_BEG2_input[1]),
    .A2(J_l_AB_BEG2_input[2]),
    .A3(J_l_AB_BEG2_input[3]),
    .S0(ConfigBits[348+0]),
    .S0N(ConfigBits_N[348+0]),
    .S1(ConfigBits[348+1]),
    .S1N(ConfigBits_N[348+1]),
    .X(J_l_AB_BEG2)
);

 //switch matrix multiplexer J_l_AB_BEG3 MUX-4
assign J_l_AB_BEG3_input = {JW2END1,S4END0,E6END0,N4END0};
cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG3 (
    .A0(J_l_AB_BEG3_input[0]),
    .A1(J_l_AB_BEG3_input[1]),
    .A2(J_l_AB_BEG3_input[2]),
    .A3(J_l_AB_BEG3_input[3]),
    .S0(ConfigBits[350+0]),
    .S0N(ConfigBits_N[350+0]),
    .S1(ConfigBits[350+1]),
    .S1N(ConfigBits_N[350+1]),
    .X(J_l_AB_BEG3)
);

 //switch matrix multiplexer J_l_CD_BEG0 MUX-4
assign J_l_CD_BEG0_input = {JN2END2,WW4END2,SS4END3,E2END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG0 (
    .A0(J_l_CD_BEG0_input[0]),
    .A1(J_l_CD_BEG0_input[1]),
    .A2(J_l_CD_BEG0_input[2]),
    .A3(J_l_CD_BEG0_input[3]),
    .S0(ConfigBits[352+0]),
    .S0N(ConfigBits_N[352+0]),
    .S1(ConfigBits[352+1]),
    .S1N(ConfigBits_N[352+1]),
    .X(J_l_CD_BEG0)
);

 //switch matrix multiplexer J_l_CD_BEG1 MUX-4
assign J_l_CD_BEG1_input = {JE2END2,W2END7,E2END2,N4END2};
cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG1 (
    .A0(J_l_CD_BEG1_input[0]),
    .A1(J_l_CD_BEG1_input[1]),
    .A2(J_l_CD_BEG1_input[2]),
    .A3(J_l_CD_BEG1_input[3]),
    .S0(ConfigBits[354+0]),
    .S0N(ConfigBits_N[354+0]),
    .S1(ConfigBits[354+1]),
    .S1N(ConfigBits_N[354+1]),
    .X(J_l_CD_BEG1)
);

 //switch matrix multiplexer J_l_CD_BEG2 MUX-4
assign J_l_CD_BEG2_input = {JS2END2,S4END1,EE4END1,NN4END1};
cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG2 (
    .A0(J_l_CD_BEG2_input[0]),
    .A1(J_l_CD_BEG2_input[1]),
    .A2(J_l_CD_BEG2_input[2]),
    .A3(J_l_CD_BEG2_input[3]),
    .S0(ConfigBits[356+0]),
    .S0N(ConfigBits_N[356+0]),
    .S1(ConfigBits[356+1]),
    .S1N(ConfigBits_N[356+1]),
    .X(J_l_CD_BEG2)
);

 //switch matrix multiplexer J_l_CD_BEG3 MUX-4
assign J_l_CD_BEG3_input = {JW2END2,W6END0,SS4END0,N4END0};
cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG3 (
    .A0(J_l_CD_BEG3_input[0]),
    .A1(J_l_CD_BEG3_input[1]),
    .A2(J_l_CD_BEG3_input[2]),
    .A3(J_l_CD_BEG3_input[3]),
    .S0(ConfigBits[358+0]),
    .S0N(ConfigBits_N[358+0]),
    .S1(ConfigBits[358+1]),
    .S1N(ConfigBits_N[358+1]),
    .X(J_l_CD_BEG3)
);

 //switch matrix multiplexer J_l_EF_BEG0 MUX-4
assign J_l_EF_BEG0_input = {JN2END3,W2END3,E2END3,N4END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG0 (
    .A0(J_l_EF_BEG0_input[0]),
    .A1(J_l_EF_BEG0_input[1]),
    .A2(J_l_EF_BEG0_input[2]),
    .A3(J_l_EF_BEG0_input[3]),
    .S0(ConfigBits[360+0]),
    .S0N(ConfigBits_N[360+0]),
    .S1(ConfigBits[360+1]),
    .S1N(ConfigBits_N[360+1]),
    .X(J_l_EF_BEG0)
);

 //switch matrix multiplexer J_l_EF_BEG1 MUX-4
assign J_l_EF_BEG1_input = {JE2END3,S4END2,E2END2,NN4END2};
cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG1 (
    .A0(J_l_EF_BEG1_input[0]),
    .A1(J_l_EF_BEG1_input[1]),
    .A2(J_l_EF_BEG1_input[2]),
    .A3(J_l_EF_BEG1_input[3]),
    .S0(ConfigBits[362+0]),
    .S0N(ConfigBits_N[362+0]),
    .S1(ConfigBits[362+1]),
    .S1N(ConfigBits_N[362+1]),
    .X(J_l_EF_BEG1)
);

 //switch matrix multiplexer J_l_EF_BEG2 MUX-4
assign J_l_EF_BEG2_input = {JS2END3,W2END4,SS4END1,N4END1};
cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG2 (
    .A0(J_l_EF_BEG2_input[0]),
    .A1(J_l_EF_BEG2_input[1]),
    .A2(J_l_EF_BEG2_input[2]),
    .A3(J_l_EF_BEG2_input[3]),
    .S0(ConfigBits[364+0]),
    .S0N(ConfigBits_N[364+0]),
    .S1(ConfigBits[364+1]),
    .S1N(ConfigBits_N[364+1]),
    .X(J_l_EF_BEG2)
);

 //switch matrix multiplexer J_l_EF_BEG3 MUX-4
assign J_l_EF_BEG3_input = {JW2END3,WW4END1,S4END0,EE4END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG3 (
    .A0(J_l_EF_BEG3_input[0]),
    .A1(J_l_EF_BEG3_input[1]),
    .A2(J_l_EF_BEG3_input[2]),
    .A3(J_l_EF_BEG3_input[3]),
    .S0(ConfigBits[366+0]),
    .S0N(ConfigBits_N[366+0]),
    .S1(ConfigBits[366+1]),
    .S1N(ConfigBits_N[366+1]),
    .X(J_l_EF_BEG3)
);

 //switch matrix multiplexer J_l_GH_BEG0 MUX-4
assign J_l_GH_BEG0_input = {JN2END4,S4END3,EE4END0,N4END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG0 (
    .A0(J_l_GH_BEG0_input[0]),
    .A1(J_l_GH_BEG0_input[1]),
    .A2(J_l_GH_BEG0_input[2]),
    .A3(J_l_GH_BEG0_input[3]),
    .S0(ConfigBits[368+0]),
    .S0N(ConfigBits_N[368+0]),
    .S1(ConfigBits[368+1]),
    .S1N(ConfigBits_N[368+1]),
    .X(J_l_GH_BEG0)
);

 //switch matrix multiplexer J_l_GH_BEG1 MUX-4
assign J_l_GH_BEG1_input = {JE2END4,W2END2,SS4END2,N4END2};
cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG1 (
    .A0(J_l_GH_BEG1_input[0]),
    .A1(J_l_GH_BEG1_input[1]),
    .A2(J_l_GH_BEG1_input[2]),
    .A3(J_l_GH_BEG1_input[3]),
    .S0(ConfigBits[370+0]),
    .S0N(ConfigBits_N[370+0]),
    .S1(ConfigBits[370+1]),
    .S1N(ConfigBits_N[370+1]),
    .X(J_l_GH_BEG1)
);

 //switch matrix multiplexer J_l_GH_BEG2 MUX-4
assign J_l_GH_BEG2_input = {JS2END4,WW4END3,S4END1,E6END1};
cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG2 (
    .A0(J_l_GH_BEG2_input[0]),
    .A1(J_l_GH_BEG2_input[1]),
    .A2(J_l_GH_BEG2_input[2]),
    .A3(J_l_GH_BEG2_input[3]),
    .S0(ConfigBits[372+0]),
    .S0N(ConfigBits_N[372+0]),
    .S1(ConfigBits[372+1]),
    .S1N(ConfigBits_N[372+1]),
    .X(J_l_GH_BEG2)
);

 //switch matrix multiplexer J_l_GH_BEG3 MUX-4
assign J_l_GH_BEG3_input = {JW2END4,W2END0,E6END0,NN4END0};
cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG3 (
    .A0(J_l_GH_BEG3_input[0]),
    .A1(J_l_GH_BEG3_input[1]),
    .A2(J_l_GH_BEG3_input[2]),
    .A3(J_l_GH_BEG3_input[3]),
    .S0(ConfigBits[374+0]),
    .S0N(ConfigBits_N[374+0]),
    .S1(ConfigBits[374+1]),
    .S1N(ConfigBits_N[374+1]),
    .X(J_l_GH_BEG3)
);


assign DEBUG_select_N1BEG0          = ConfigBits[1:0];
assign DEBUG_select_N1BEG1          = ConfigBits[3:2];
assign DEBUG_select_N1BEG2          = ConfigBits[5:4];
assign DEBUG_select_N1BEG3          = ConfigBits[7:6];
assign DEBUG_select_N4BEG0          = ConfigBits[9:8];
assign DEBUG_select_N4BEG1          = ConfigBits[11:10];
assign DEBUG_select_N4BEG2          = ConfigBits[13:12];
assign DEBUG_select_N4BEG3          = ConfigBits[15:14];
assign DEBUG_select_NN4BEG0         = ConfigBits[18:16];
assign DEBUG_select_NN4BEG1         = ConfigBits[21:19];
assign DEBUG_select_NN4BEG2         = ConfigBits[24:22];
assign DEBUG_select_NN4BEG3         = ConfigBits[27:25];
assign DEBUG_select_E1BEG0          = ConfigBits[29:28];
assign DEBUG_select_E1BEG1          = ConfigBits[31:30];
assign DEBUG_select_E1BEG2          = ConfigBits[33:32];
assign DEBUG_select_E1BEG3          = ConfigBits[35:34];
assign DEBUG_select_EE4BEG0         = ConfigBits[38:36];
assign DEBUG_select_EE4BEG1         = ConfigBits[41:39];
assign DEBUG_select_EE4BEG2         = ConfigBits[44:42];
assign DEBUG_select_EE4BEG3         = ConfigBits[47:45];
assign DEBUG_select_E6BEG0          = ConfigBits[51:48];
assign DEBUG_select_E6BEG1          = ConfigBits[55:52];
assign DEBUG_select_S1BEG0          = ConfigBits[57:56];
assign DEBUG_select_S1BEG1          = ConfigBits[59:58];
assign DEBUG_select_S1BEG2          = ConfigBits[61:60];
assign DEBUG_select_S1BEG3          = ConfigBits[63:62];
assign DEBUG_select_S4BEG0          = ConfigBits[65:64];
assign DEBUG_select_S4BEG1          = ConfigBits[67:66];
assign DEBUG_select_S4BEG2          = ConfigBits[69:68];
assign DEBUG_select_S4BEG3          = ConfigBits[71:70];
assign DEBUG_select_SS4BEG0         = ConfigBits[74:72];
assign DEBUG_select_SS4BEG1         = ConfigBits[77:75];
assign DEBUG_select_SS4BEG2         = ConfigBits[80:78];
assign DEBUG_select_SS4BEG3         = ConfigBits[83:81];
assign DEBUG_select_W1BEG0          = ConfigBits[85:84];
assign DEBUG_select_W1BEG1          = ConfigBits[87:86];
assign DEBUG_select_W1BEG2          = ConfigBits[89:88];
assign DEBUG_select_W1BEG3          = ConfigBits[91:90];
assign DEBUG_select_WW4BEG0         = ConfigBits[94:92];
assign DEBUG_select_WW4BEG1         = ConfigBits[97:95];
assign DEBUG_select_WW4BEG2         = ConfigBits[100:98];
assign DEBUG_select_WW4BEG3         = ConfigBits[103:101];
assign DEBUG_select_W6BEG0          = ConfigBits[107:104];
assign DEBUG_select_W6BEG1          = ConfigBits[111:108];
assign DEBUG_select_resp_ready      = ConfigBits[113:112];
assign DEBUG_select_t_req_ready     = ConfigBits[115:114];
assign DEBUG_select_t_resp_status0  = ConfigBits[117:116];
assign DEBUG_select_t_resp_status1  = ConfigBits[119:118];
assign DEBUG_select_t_resp_status2  = ConfigBits[121:120];
assign DEBUG_select_t_resp_valid    = ConfigBits[123:122];
assign DEBUG_select_J2MID_ABa_BEG0  = ConfigBits[125:124];
assign DEBUG_select_J2MID_ABa_BEG1  = ConfigBits[127:126];
assign DEBUG_select_J2MID_ABa_BEG2  = ConfigBits[129:128];
assign DEBUG_select_J2MID_ABa_BEG3  = ConfigBits[131:130];
assign DEBUG_select_J2MID_CDa_BEG0  = ConfigBits[133:132];
assign DEBUG_select_J2MID_CDa_BEG1  = ConfigBits[135:134];
assign DEBUG_select_J2MID_CDa_BEG2  = ConfigBits[137:136];
assign DEBUG_select_J2MID_CDa_BEG3  = ConfigBits[139:138];
assign DEBUG_select_J2MID_EFa_BEG0  = ConfigBits[141:140];
assign DEBUG_select_J2MID_EFa_BEG1  = ConfigBits[143:142];
assign DEBUG_select_J2MID_EFa_BEG2  = ConfigBits[145:144];
assign DEBUG_select_J2MID_EFa_BEG3  = ConfigBits[147:146];
assign DEBUG_select_J2MID_GHa_BEG0  = ConfigBits[149:148];
assign DEBUG_select_J2MID_GHa_BEG1  = ConfigBits[151:150];
assign DEBUG_select_J2MID_GHa_BEG2  = ConfigBits[153:152];
assign DEBUG_select_J2MID_GHa_BEG3  = ConfigBits[155:154];
assign DEBUG_select_J2MID_ABb_BEG0  = ConfigBits[157:156];
assign DEBUG_select_J2MID_ABb_BEG1  = ConfigBits[159:158];
assign DEBUG_select_J2MID_ABb_BEG2  = ConfigBits[161:160];
assign DEBUG_select_J2MID_ABb_BEG3  = ConfigBits[163:162];
assign DEBUG_select_J2MID_CDb_BEG0  = ConfigBits[165:164];
assign DEBUG_select_J2MID_CDb_BEG1  = ConfigBits[167:166];
assign DEBUG_select_J2MID_CDb_BEG2  = ConfigBits[169:168];
assign DEBUG_select_J2MID_CDb_BEG3  = ConfigBits[171:170];
assign DEBUG_select_J2MID_EFb_BEG0  = ConfigBits[173:172];
assign DEBUG_select_J2MID_EFb_BEG1  = ConfigBits[175:174];
assign DEBUG_select_J2MID_EFb_BEG2  = ConfigBits[177:176];
assign DEBUG_select_J2MID_EFb_BEG3  = ConfigBits[179:178];
assign DEBUG_select_J2MID_GHb_BEG0  = ConfigBits[181:180];
assign DEBUG_select_J2MID_GHb_BEG1  = ConfigBits[183:182];
assign DEBUG_select_J2MID_GHb_BEG2  = ConfigBits[185:184];
assign DEBUG_select_J2MID_GHb_BEG3  = ConfigBits[187:186];
assign DEBUG_select_J2END_AB_BEG0   = ConfigBits[189:188];
assign DEBUG_select_J2END_AB_BEG1   = ConfigBits[191:190];
assign DEBUG_select_J2END_AB_BEG2   = ConfigBits[193:192];
assign DEBUG_select_J2END_AB_BEG3   = ConfigBits[195:194];
assign DEBUG_select_J2END_CD_BEG0   = ConfigBits[197:196];
assign DEBUG_select_J2END_CD_BEG1   = ConfigBits[199:198];
assign DEBUG_select_J2END_CD_BEG2   = ConfigBits[201:200];
assign DEBUG_select_J2END_CD_BEG3   = ConfigBits[203:202];
assign DEBUG_select_J2END_EF_BEG0   = ConfigBits[205:204];
assign DEBUG_select_J2END_EF_BEG1   = ConfigBits[207:206];
assign DEBUG_select_J2END_EF_BEG2   = ConfigBits[209:208];
assign DEBUG_select_J2END_EF_BEG3   = ConfigBits[211:210];
assign DEBUG_select_J2END_GH_BEG0   = ConfigBits[213:212];
assign DEBUG_select_J2END_GH_BEG1   = ConfigBits[215:214];
assign DEBUG_select_J2END_GH_BEG2   = ConfigBits[217:216];
assign DEBUG_select_J2END_GH_BEG3   = ConfigBits[219:218];
assign DEBUG_select_JN2BEG0         = ConfigBits[223:220];
assign DEBUG_select_JN2BEG1         = ConfigBits[227:224];
assign DEBUG_select_JN2BEG2         = ConfigBits[231:228];
assign DEBUG_select_JN2BEG3         = ConfigBits[235:232];
assign DEBUG_select_JN2BEG4         = ConfigBits[239:236];
assign DEBUG_select_JN2BEG5         = ConfigBits[243:240];
assign DEBUG_select_JN2BEG6         = ConfigBits[247:244];
assign DEBUG_select_JN2BEG7         = ConfigBits[251:248];
assign DEBUG_select_JE2BEG0         = ConfigBits[255:252];
assign DEBUG_select_JE2BEG1         = ConfigBits[259:256];
assign DEBUG_select_JE2BEG2         = ConfigBits[263:260];
assign DEBUG_select_JE2BEG3         = ConfigBits[267:264];
assign DEBUG_select_JE2BEG4         = ConfigBits[271:268];
assign DEBUG_select_JE2BEG5         = ConfigBits[275:272];
assign DEBUG_select_JE2BEG6         = ConfigBits[279:276];
assign DEBUG_select_JE2BEG7         = ConfigBits[283:280];
assign DEBUG_select_JS2BEG0         = ConfigBits[287:284];
assign DEBUG_select_JS2BEG1         = ConfigBits[291:288];
assign DEBUG_select_JS2BEG2         = ConfigBits[295:292];
assign DEBUG_select_JS2BEG3         = ConfigBits[299:296];
assign DEBUG_select_JS2BEG4         = ConfigBits[303:300];
assign DEBUG_select_JS2BEG5         = ConfigBits[307:304];
assign DEBUG_select_JS2BEG6         = ConfigBits[311:308];
assign DEBUG_select_JS2BEG7         = ConfigBits[315:312];
assign DEBUG_select_JW2BEG0         = ConfigBits[319:316];
assign DEBUG_select_JW2BEG1         = ConfigBits[323:320];
assign DEBUG_select_JW2BEG2         = ConfigBits[327:324];
assign DEBUG_select_JW2BEG3         = ConfigBits[331:328];
assign DEBUG_select_JW2BEG4         = ConfigBits[335:332];
assign DEBUG_select_JW2BEG5         = ConfigBits[339:336];
assign DEBUG_select_JW2BEG6         = ConfigBits[343:340];
assign DEBUG_select_JW2BEG7         = ConfigBits[347:344];
assign DEBUG_select_J_l_AB_BEG0     = ConfigBits[349:348];
assign DEBUG_select_J_l_AB_BEG1     = ConfigBits[351:350];
assign DEBUG_select_J_l_AB_BEG2     = ConfigBits[353:352];
assign DEBUG_select_J_l_AB_BEG3     = ConfigBits[355:354];
assign DEBUG_select_J_l_CD_BEG0     = ConfigBits[357:356];
assign DEBUG_select_J_l_CD_BEG1     = ConfigBits[359:358];
assign DEBUG_select_J_l_CD_BEG2     = ConfigBits[361:360];
assign DEBUG_select_J_l_CD_BEG3     = ConfigBits[363:362];
assign DEBUG_select_J_l_EF_BEG0     = ConfigBits[365:364];
assign DEBUG_select_J_l_EF_BEG1     = ConfigBits[367:366];
assign DEBUG_select_J_l_EF_BEG2     = ConfigBits[369:368];
assign DEBUG_select_J_l_EF_BEG3     = ConfigBits[371:370];
assign DEBUG_select_J_l_GH_BEG0     = ConfigBits[373:372];
assign DEBUG_select_J_l_GH_BEG1     = ConfigBits[375:374];
assign DEBUG_select_J_l_GH_BEG2     = ConfigBits[377:376];
assign DEBUG_select_J_l_GH_BEG3     = ConfigBits[379:378];
endmodule