 // NumberOfConfigBits: 360
module SCC2_switch_matrix
    #(
        parameter NoConfigBits=360
    )
    (
        input o_6to20,
        input o_6to21,
        input o_6to22,
        input o_6to23,
        input o_6to24,
        input o_6to25,
        input o_6to26,
        input o_6to27,
        input o_6to28,
        input o_6to29,
        input o_6to210,
        input o_6to211,
        input o_6to212,
        input o_6to213,
        input o_6to214,
        input o_6to215,
        input o_6to216,
        input o_6to217,
        input o_6to218,
        input o_6to219,
        input o_6to220,
        input o_6to221,
        input o_6to222,
        input o_6to223,
        input o_6to224,
        input o_6to225,
        input o_6to226,
        input o_6to227,
        input o_6to228,
        input o_6to229,
        input o_6to230,
        input o_6to231,
        input N1END0,
        input N1END1,
        input N1END2,
        input N1END3,
        input N2MID0,
        input N2MID1,
        input N2MID2,
        input N2MID3,
        input N2MID4,
        input N2MID5,
        input N2MID6,
        input N2MID7,
        input N2END0,
        input N2END1,
        input N2END2,
        input N2END3,
        input N2END4,
        input N2END5,
        input N2END6,
        input N2END7,
        input N4END0,
        input N4END1,
        input N4END2,
        input N4END3,
        input NN4END0,
        input NN4END1,
        input NN4END2,
        input NN4END3,
        input E1END0,
        input E1END1,
        input E1END2,
        input E1END3,
        input E2MID0,
        input E2MID1,
        input E2MID2,
        input E2MID3,
        input E2MID4,
        input E2MID5,
        input E2MID6,
        input E2MID7,
        input E2END0,
        input E2END1,
        input E2END2,
        input E2END3,
        input E2END4,
        input E2END5,
        input E2END6,
        input E2END7,
        input EE4END0,
        input EE4END1,
        input EE4END2,
        input EE4END3,
        input E6END0,
        input E6END1,
        input S1END0,
        input S1END1,
        input S1END2,
        input S1END3,
        input S2MID0,
        input S2MID1,
        input S2MID2,
        input S2MID3,
        input S2MID4,
        input S2MID5,
        input S2MID6,
        input S2MID7,
        input S2END0,
        input S2END1,
        input S2END2,
        input S2END3,
        input S2END4,
        input S2END5,
        input S2END6,
        input S2END7,
        input S4END0,
        input S4END1,
        input S4END2,
        input S4END3,
        input SS4END0,
        input SS4END1,
        input SS4END2,
        input SS4END3,
        input W1END0,
        input W1END1,
        input W1END2,
        input W1END3,
        input W2MID0,
        input W2MID1,
        input W2MID2,
        input W2MID3,
        input W2MID4,
        input W2MID5,
        input W2MID6,
        input W2MID7,
        input W2END0,
        input W2END1,
        input W2END2,
        input W2END3,
        input W2END4,
        input W2END5,
        input W2END6,
        input W2END7,
        input WW4END0,
        input WW4END1,
        input WW4END2,
        input WW4END3,
        input W6END0,
        input W6END1,
        input J2MID_ABa_END0,
        input J2MID_ABa_END1,
        input J2MID_ABa_END2,
        input J2MID_ABa_END3,
        input J2MID_CDa_END0,
        input J2MID_CDa_END1,
        input J2MID_CDa_END2,
        input J2MID_CDa_END3,
        input J2MID_EFa_END0,
        input J2MID_EFa_END1,
        input J2MID_EFa_END2,
        input J2MID_EFa_END3,
        input J2MID_GHa_END0,
        input J2MID_GHa_END1,
        input J2MID_GHa_END2,
        input J2MID_GHa_END3,
        input J2MID_ABb_END0,
        input J2MID_ABb_END1,
        input J2MID_ABb_END2,
        input J2MID_ABb_END3,
        input J2MID_CDb_END0,
        input J2MID_CDb_END1,
        input J2MID_CDb_END2,
        input J2MID_CDb_END3,
        input J2MID_EFb_END0,
        input J2MID_EFb_END1,
        input J2MID_EFb_END2,
        input J2MID_EFb_END3,
        input J2MID_GHb_END0,
        input J2MID_GHb_END1,
        input J2MID_GHb_END2,
        input J2MID_GHb_END3,
        input J2END_AB_END0,
        input J2END_AB_END1,
        input J2END_AB_END2,
        input J2END_AB_END3,
        input J2END_CD_END0,
        input J2END_CD_END1,
        input J2END_CD_END2,
        input J2END_CD_END3,
        input J2END_EF_END0,
        input J2END_EF_END1,
        input J2END_EF_END2,
        input J2END_EF_END3,
        input J2END_GH_END0,
        input J2END_GH_END1,
        input J2END_GH_END2,
        input J2END_GH_END3,
        input JN2END0,
        input JN2END1,
        input JN2END2,
        input JN2END3,
        input JN2END4,
        input JN2END5,
        input JN2END6,
        input JN2END7,
        input JE2END0,
        input JE2END1,
        input JE2END2,
        input JE2END3,
        input JE2END4,
        input JE2END5,
        input JE2END6,
        input JE2END7,
        input JS2END0,
        input JS2END1,
        input JS2END2,
        input JS2END3,
        input JS2END4,
        input JS2END5,
        input JS2END6,
        input JS2END7,
        input JW2END0,
        input JW2END1,
        input JW2END2,
        input JW2END3,
        input JW2END4,
        input JW2END5,
        input JW2END6,
        input JW2END7,
        input J_l_AB_END0,
        input J_l_AB_END1,
        input J_l_AB_END2,
        input J_l_AB_END3,
        input J_l_CD_END0,
        input J_l_CD_END1,
        input J_l_CD_END2,
        input J_l_CD_END3,
        input J_l_EF_END0,
        input J_l_EF_END1,
        input J_l_EF_END2,
        input J_l_EF_END3,
        input J_l_GH_END0,
        input J_l_GH_END1,
        input J_l_GH_END2,
        input J_l_GH_END3,
        output i_2to60,
        output i_2to61,
        output i_2to62,
        output i_2to63,
        output i_2to64,
        output i_2to65,
        output i_2to66,
        output i_2to67,
        output i_2to68,
        output i_2to69,
        output i_2to610,
        output i_2to611,
        output i_2to612,
        output i_2to613,
        output i_2to614,
        output i_2to615,
        output i_2to616,
        output i_2to617,
        output i_2to618,
        output i_2to619,
        output i_2to620,
        output i_2to621,
        output i_2to622,
        output i_2to623,
        output i_2to624,
        output i_2to625,
        output i_2to626,
        output i_2to627,
        output i_2to628,
        output i_2to629,
        output i_2to630,
        output i_2to631,
        output N1BEG0,
        output N1BEG1,
        output N1BEG2,
        output N1BEG3,
        output N2BEG0,
        output N2BEG1,
        output N2BEG2,
        output N2BEG3,
        output N2BEG4,
        output N2BEG5,
        output N2BEG6,
        output N2BEG7,
        output N2BEGb0,
        output N2BEGb1,
        output N2BEGb2,
        output N2BEGb3,
        output N2BEGb4,
        output N2BEGb5,
        output N2BEGb6,
        output N2BEGb7,
        output N4BEG0,
        output N4BEG1,
        output N4BEG2,
        output N4BEG3,
        output NN4BEG0,
        output NN4BEG1,
        output NN4BEG2,
        output NN4BEG3,
        output E1BEG0,
        output E1BEG1,
        output E1BEG2,
        output E1BEG3,
        output E2BEG0,
        output E2BEG1,
        output E2BEG2,
        output E2BEG3,
        output E2BEG4,
        output E2BEG5,
        output E2BEG6,
        output E2BEG7,
        output E2BEGb0,
        output E2BEGb1,
        output E2BEGb2,
        output E2BEGb3,
        output E2BEGb4,
        output E2BEGb5,
        output E2BEGb6,
        output E2BEGb7,
        output EE4BEG0,
        output EE4BEG1,
        output EE4BEG2,
        output EE4BEG3,
        output E6BEG0,
        output E6BEG1,
        output S1BEG0,
        output S1BEG1,
        output S1BEG2,
        output S1BEG3,
        output S2BEG0,
        output S2BEG1,
        output S2BEG2,
        output S2BEG3,
        output S2BEG4,
        output S2BEG5,
        output S2BEG6,
        output S2BEG7,
        output S2BEGb0,
        output S2BEGb1,
        output S2BEGb2,
        output S2BEGb3,
        output S2BEGb4,
        output S2BEGb5,
        output S2BEGb6,
        output S2BEGb7,
        output S4BEG0,
        output S4BEG1,
        output S4BEG2,
        output S4BEG3,
        output SS4BEG0,
        output SS4BEG1,
        output SS4BEG2,
        output SS4BEG3,
        output W1BEG0,
        output W1BEG1,
        output W1BEG2,
        output W1BEG3,
        output W2BEG0,
        output W2BEG1,
        output W2BEG2,
        output W2BEG3,
        output W2BEG4,
        output W2BEG5,
        output W2BEG6,
        output W2BEG7,
        output W2BEGb0,
        output W2BEGb1,
        output W2BEGb2,
        output W2BEGb3,
        output W2BEGb4,
        output W2BEGb5,
        output W2BEGb6,
        output W2BEGb7,
        output WW4BEG0,
        output WW4BEG1,
        output WW4BEG2,
        output WW4BEG3,
        output W6BEG0,
        output W6BEG1,
        output J2MID_ABa_BEG0,
        output J2MID_ABa_BEG1,
        output J2MID_ABa_BEG2,
        output J2MID_ABa_BEG3,
        output J2MID_CDa_BEG0,
        output J2MID_CDa_BEG1,
        output J2MID_CDa_BEG2,
        output J2MID_CDa_BEG3,
        output J2MID_EFa_BEG0,
        output J2MID_EFa_BEG1,
        output J2MID_EFa_BEG2,
        output J2MID_EFa_BEG3,
        output J2MID_GHa_BEG0,
        output J2MID_GHa_BEG1,
        output J2MID_GHa_BEG2,
        output J2MID_GHa_BEG3,
        output J2MID_ABb_BEG0,
        output J2MID_ABb_BEG1,
        output J2MID_ABb_BEG2,
        output J2MID_ABb_BEG3,
        output J2MID_CDb_BEG0,
        output J2MID_CDb_BEG1,
        output J2MID_CDb_BEG2,
        output J2MID_CDb_BEG3,
        output J2MID_EFb_BEG0,
        output J2MID_EFb_BEG1,
        output J2MID_EFb_BEG2,
        output J2MID_EFb_BEG3,
        output J2MID_GHb_BEG0,
        output J2MID_GHb_BEG1,
        output J2MID_GHb_BEG2,
        output J2MID_GHb_BEG3,
        output J2END_AB_BEG0,
        output J2END_AB_BEG1,
        output J2END_AB_BEG2,
        output J2END_AB_BEG3,
        output J2END_CD_BEG0,
        output J2END_CD_BEG1,
        output J2END_CD_BEG2,
        output J2END_CD_BEG3,
        output J2END_EF_BEG0,
        output J2END_EF_BEG1,
        output J2END_EF_BEG2,
        output J2END_EF_BEG3,
        output J2END_GH_BEG0,
        output J2END_GH_BEG1,
        output J2END_GH_BEG2,
        output J2END_GH_BEG3,
        output JN2BEG0,
        output JN2BEG1,
        output JN2BEG2,
        output JN2BEG3,
        output JN2BEG4,
        output JN2BEG5,
        output JN2BEG6,
        output JN2BEG7,
        output JE2BEG0,
        output JE2BEG1,
        output JE2BEG2,
        output JE2BEG3,
        output JE2BEG4,
        output JE2BEG5,
        output JE2BEG6,
        output JE2BEG7,
        output JS2BEG0,
        output JS2BEG1,
        output JS2BEG2,
        output JS2BEG3,
        output JS2BEG4,
        output JS2BEG5,
        output JS2BEG6,
        output JS2BEG7,
        output JW2BEG0,
        output JW2BEG1,
        output JW2BEG2,
        output JW2BEG3,
        output JW2BEG4,
        output JW2BEG5,
        output JW2BEG6,
        output JW2BEG7,
        output J_l_AB_BEG0,
        output J_l_AB_BEG1,
        output J_l_AB_BEG2,
        output J_l_AB_BEG3,
        output J_l_CD_BEG0,
        output J_l_CD_BEG1,
        output J_l_CD_BEG2,
        output J_l_CD_BEG3,
        output J_l_EF_BEG0,
        output J_l_EF_BEG1,
        output J_l_EF_BEG2,
        output J_l_EF_BEG3,
        output J_l_GH_BEG0,
        output J_l_GH_BEG1,
        output J_l_GH_BEG2,
        output J_l_GH_BEG3,
 //global
        input [NoConfigBits-1:0] ConfigBits,
        input [NoConfigBits-1:0] ConfigBits_N
);
parameter GND0 = 1'b0;
parameter GND = 1'b0;
parameter VCC0 = 1'b1;
parameter VCC = 1'b1;
parameter VDD0 = 1'b1;
parameter VDD = 1'b1;

wire[4-1:0] i_2to60_input;
wire[4-1:0] i_2to61_input;
wire[4-1:0] i_2to62_input;
wire[4-1:0] i_2to63_input;
wire[4-1:0] i_2to64_input;
wire[4-1:0] i_2to65_input;
wire[4-1:0] i_2to66_input;
wire[4-1:0] i_2to67_input;
wire[0-1:0] i_2to68_input;
wire[0-1:0] i_2to69_input;
wire[0-1:0] i_2to610_input;
wire[0-1:0] i_2to611_input;
wire[0-1:0] i_2to612_input;
wire[0-1:0] i_2to613_input;
wire[0-1:0] i_2to614_input;
wire[0-1:0] i_2to615_input;
wire[0-1:0] i_2to616_input;
wire[0-1:0] i_2to617_input;
wire[0-1:0] i_2to618_input;
wire[0-1:0] i_2to619_input;
wire[0-1:0] i_2to620_input;
wire[0-1:0] i_2to621_input;
wire[0-1:0] i_2to622_input;
wire[0-1:0] i_2to623_input;
wire[0-1:0] i_2to624_input;
wire[0-1:0] i_2to625_input;
wire[0-1:0] i_2to626_input;
wire[0-1:0] i_2to627_input;
wire[0-1:0] i_2to628_input;
wire[0-1:0] i_2to629_input;
wire[0-1:0] i_2to630_input;
wire[0-1:0] i_2to631_input;
wire[4-1:0] N1BEG0_input;
wire[4-1:0] N1BEG1_input;
wire[4-1:0] N1BEG2_input;
wire[4-1:0] N1BEG3_input;
wire[1-1:0] N2BEG0_input;
wire[1-1:0] N2BEG1_input;
wire[1-1:0] N2BEG2_input;
wire[1-1:0] N2BEG3_input;
wire[1-1:0] N2BEG4_input;
wire[1-1:0] N2BEG5_input;
wire[1-1:0] N2BEG6_input;
wire[1-1:0] N2BEG7_input;
wire[1-1:0] N2BEGb0_input;
wire[1-1:0] N2BEGb1_input;
wire[1-1:0] N2BEGb2_input;
wire[1-1:0] N2BEGb3_input;
wire[1-1:0] N2BEGb4_input;
wire[1-1:0] N2BEGb5_input;
wire[1-1:0] N2BEGb6_input;
wire[1-1:0] N2BEGb7_input;
wire[4-1:0] N4BEG0_input;
wire[4-1:0] N4BEG1_input;
wire[4-1:0] N4BEG2_input;
wire[4-1:0] N4BEG3_input;
wire[8-1:0] NN4BEG0_input;
wire[8-1:0] NN4BEG1_input;
wire[8-1:0] NN4BEG2_input;
wire[8-1:0] NN4BEG3_input;
wire[4-1:0] E1BEG0_input;
wire[4-1:0] E1BEG1_input;
wire[4-1:0] E1BEG2_input;
wire[4-1:0] E1BEG3_input;
wire[1-1:0] E2BEG0_input;
wire[1-1:0] E2BEG1_input;
wire[1-1:0] E2BEG2_input;
wire[1-1:0] E2BEG3_input;
wire[1-1:0] E2BEG4_input;
wire[1-1:0] E2BEG5_input;
wire[1-1:0] E2BEG6_input;
wire[1-1:0] E2BEG7_input;
wire[1-1:0] E2BEGb0_input;
wire[1-1:0] E2BEGb1_input;
wire[1-1:0] E2BEGb2_input;
wire[1-1:0] E2BEGb3_input;
wire[1-1:0] E2BEGb4_input;
wire[1-1:0] E2BEGb5_input;
wire[1-1:0] E2BEGb6_input;
wire[1-1:0] E2BEGb7_input;
wire[8-1:0] EE4BEG0_input;
wire[8-1:0] EE4BEG1_input;
wire[8-1:0] EE4BEG2_input;
wire[8-1:0] EE4BEG3_input;
wire[16-1:0] E6BEG0_input;
wire[16-1:0] E6BEG1_input;
wire[4-1:0] S1BEG0_input;
wire[4-1:0] S1BEG1_input;
wire[4-1:0] S1BEG2_input;
wire[4-1:0] S1BEG3_input;
wire[1-1:0] S2BEG0_input;
wire[1-1:0] S2BEG1_input;
wire[1-1:0] S2BEG2_input;
wire[1-1:0] S2BEG3_input;
wire[1-1:0] S2BEG4_input;
wire[1-1:0] S2BEG5_input;
wire[1-1:0] S2BEG6_input;
wire[1-1:0] S2BEG7_input;
wire[1-1:0] S2BEGb0_input;
wire[1-1:0] S2BEGb1_input;
wire[1-1:0] S2BEGb2_input;
wire[1-1:0] S2BEGb3_input;
wire[1-1:0] S2BEGb4_input;
wire[1-1:0] S2BEGb5_input;
wire[1-1:0] S2BEGb6_input;
wire[1-1:0] S2BEGb7_input;
wire[4-1:0] S4BEG0_input;
wire[4-1:0] S4BEG1_input;
wire[4-1:0] S4BEG2_input;
wire[4-1:0] S4BEG3_input;
wire[8-1:0] SS4BEG0_input;
wire[8-1:0] SS4BEG1_input;
wire[8-1:0] SS4BEG2_input;
wire[8-1:0] SS4BEG3_input;
wire[4-1:0] W1BEG0_input;
wire[4-1:0] W1BEG1_input;
wire[4-1:0] W1BEG2_input;
wire[4-1:0] W1BEG3_input;
wire[1-1:0] W2BEG0_input;
wire[1-1:0] W2BEG1_input;
wire[1-1:0] W2BEG2_input;
wire[1-1:0] W2BEG3_input;
wire[1-1:0] W2BEG4_input;
wire[1-1:0] W2BEG5_input;
wire[1-1:0] W2BEG6_input;
wire[1-1:0] W2BEG7_input;
wire[1-1:0] W2BEGb0_input;
wire[1-1:0] W2BEGb1_input;
wire[1-1:0] W2BEGb2_input;
wire[1-1:0] W2BEGb3_input;
wire[1-1:0] W2BEGb4_input;
wire[1-1:0] W2BEGb5_input;
wire[1-1:0] W2BEGb6_input;
wire[1-1:0] W2BEGb7_input;
wire[8-1:0] WW4BEG0_input;
wire[8-1:0] WW4BEG1_input;
wire[8-1:0] WW4BEG2_input;
wire[8-1:0] WW4BEG3_input;
wire[16-1:0] W6BEG0_input;
wire[16-1:0] W6BEG1_input;
wire[4-1:0] J2MID_ABa_BEG0_input;
wire[4-1:0] J2MID_ABa_BEG1_input;
wire[4-1:0] J2MID_ABa_BEG2_input;
wire[4-1:0] J2MID_ABa_BEG3_input;
wire[4-1:0] J2MID_CDa_BEG0_input;
wire[4-1:0] J2MID_CDa_BEG1_input;
wire[4-1:0] J2MID_CDa_BEG2_input;
wire[4-1:0] J2MID_CDa_BEG3_input;
wire[4-1:0] J2MID_EFa_BEG0_input;
wire[4-1:0] J2MID_EFa_BEG1_input;
wire[4-1:0] J2MID_EFa_BEG2_input;
wire[4-1:0] J2MID_EFa_BEG3_input;
wire[4-1:0] J2MID_GHa_BEG0_input;
wire[4-1:0] J2MID_GHa_BEG1_input;
wire[4-1:0] J2MID_GHa_BEG2_input;
wire[4-1:0] J2MID_GHa_BEG3_input;
wire[4-1:0] J2MID_ABb_BEG0_input;
wire[4-1:0] J2MID_ABb_BEG1_input;
wire[4-1:0] J2MID_ABb_BEG2_input;
wire[4-1:0] J2MID_ABb_BEG3_input;
wire[4-1:0] J2MID_CDb_BEG0_input;
wire[4-1:0] J2MID_CDb_BEG1_input;
wire[4-1:0] J2MID_CDb_BEG2_input;
wire[4-1:0] J2MID_CDb_BEG3_input;
wire[4-1:0] J2MID_EFb_BEG0_input;
wire[4-1:0] J2MID_EFb_BEG1_input;
wire[4-1:0] J2MID_EFb_BEG2_input;
wire[4-1:0] J2MID_EFb_BEG3_input;
wire[4-1:0] J2MID_GHb_BEG0_input;
wire[4-1:0] J2MID_GHb_BEG1_input;
wire[4-1:0] J2MID_GHb_BEG2_input;
wire[4-1:0] J2MID_GHb_BEG3_input;
wire[4-1:0] J2END_AB_BEG0_input;
wire[4-1:0] J2END_AB_BEG1_input;
wire[4-1:0] J2END_AB_BEG2_input;
wire[4-1:0] J2END_AB_BEG3_input;
wire[4-1:0] J2END_CD_BEG0_input;
wire[4-1:0] J2END_CD_BEG1_input;
wire[4-1:0] J2END_CD_BEG2_input;
wire[4-1:0] J2END_CD_BEG3_input;
wire[4-1:0] J2END_EF_BEG0_input;
wire[4-1:0] J2END_EF_BEG1_input;
wire[4-1:0] J2END_EF_BEG2_input;
wire[4-1:0] J2END_EF_BEG3_input;
wire[4-1:0] J2END_GH_BEG0_input;
wire[4-1:0] J2END_GH_BEG1_input;
wire[4-1:0] J2END_GH_BEG2_input;
wire[4-1:0] J2END_GH_BEG3_input;
wire[16-1:0] JN2BEG0_input;
wire[16-1:0] JN2BEG1_input;
wire[16-1:0] JN2BEG2_input;
wire[16-1:0] JN2BEG3_input;
wire[16-1:0] JN2BEG4_input;
wire[16-1:0] JN2BEG5_input;
wire[16-1:0] JN2BEG6_input;
wire[16-1:0] JN2BEG7_input;
wire[16-1:0] JE2BEG0_input;
wire[16-1:0] JE2BEG1_input;
wire[16-1:0] JE2BEG2_input;
wire[16-1:0] JE2BEG3_input;
wire[16-1:0] JE2BEG4_input;
wire[16-1:0] JE2BEG5_input;
wire[16-1:0] JE2BEG6_input;
wire[16-1:0] JE2BEG7_input;
wire[16-1:0] JS2BEG0_input;
wire[16-1:0] JS2BEG1_input;
wire[16-1:0] JS2BEG2_input;
wire[16-1:0] JS2BEG3_input;
wire[16-1:0] JS2BEG4_input;
wire[16-1:0] JS2BEG5_input;
wire[16-1:0] JS2BEG6_input;
wire[16-1:0] JS2BEG7_input;
wire[16-1:0] JW2BEG0_input;
wire[16-1:0] JW2BEG1_input;
wire[16-1:0] JW2BEG2_input;
wire[16-1:0] JW2BEG3_input;
wire[16-1:0] JW2BEG4_input;
wire[16-1:0] JW2BEG5_input;
wire[16-1:0] JW2BEG6_input;
wire[16-1:0] JW2BEG7_input;
wire[4-1:0] J_l_AB_BEG0_input;
wire[4-1:0] J_l_AB_BEG1_input;
wire[4-1:0] J_l_AB_BEG2_input;
wire[4-1:0] J_l_AB_BEG3_input;
wire[4-1:0] J_l_CD_BEG0_input;
wire[4-1:0] J_l_CD_BEG1_input;
wire[4-1:0] J_l_CD_BEG2_input;
wire[4-1:0] J_l_CD_BEG3_input;
wire[4-1:0] J_l_EF_BEG0_input;
wire[4-1:0] J_l_EF_BEG1_input;
wire[4-1:0] J_l_EF_BEG2_input;
wire[4-1:0] J_l_EF_BEG3_input;
wire[4-1:0] J_l_GH_BEG0_input;
wire[4-1:0] J_l_GH_BEG1_input;
wire[4-1:0] J_l_GH_BEG2_input;
wire[4-1:0] J_l_GH_BEG3_input;

wire[2-1:0] DEBUG_select_i_2to60;
wire[2-1:0] DEBUG_select_i_2to61;
wire[2-1:0] DEBUG_select_i_2to62;
wire[2-1:0] DEBUG_select_i_2to63;
wire[2-1:0] DEBUG_select_i_2to64;
wire[2-1:0] DEBUG_select_i_2to65;
wire[2-1:0] DEBUG_select_i_2to66;
wire[2-1:0] DEBUG_select_i_2to67;
wire[2-1:0] DEBUG_select_N1BEG0;
wire[2-1:0] DEBUG_select_N1BEG1;
wire[2-1:0] DEBUG_select_N1BEG2;
wire[2-1:0] DEBUG_select_N1BEG3;
wire[2-1:0] DEBUG_select_N4BEG0;
wire[2-1:0] DEBUG_select_N4BEG1;
wire[2-1:0] DEBUG_select_N4BEG2;
wire[2-1:0] DEBUG_select_N4BEG3;
wire[3-1:0] DEBUG_select_NN4BEG0;
wire[3-1:0] DEBUG_select_NN4BEG1;
wire[3-1:0] DEBUG_select_NN4BEG2;
wire[3-1:0] DEBUG_select_NN4BEG3;
wire[2-1:0] DEBUG_select_E1BEG0;
wire[2-1:0] DEBUG_select_E1BEG1;
wire[2-1:0] DEBUG_select_E1BEG2;
wire[2-1:0] DEBUG_select_E1BEG3;
wire[3-1:0] DEBUG_select_EE4BEG0;
wire[3-1:0] DEBUG_select_EE4BEG1;
wire[3-1:0] DEBUG_select_EE4BEG2;
wire[3-1:0] DEBUG_select_EE4BEG3;
wire[4-1:0] DEBUG_select_E6BEG0;
wire[4-1:0] DEBUG_select_E6BEG1;
wire[2-1:0] DEBUG_select_S1BEG0;
wire[2-1:0] DEBUG_select_S1BEG1;
wire[2-1:0] DEBUG_select_S1BEG2;
wire[2-1:0] DEBUG_select_S1BEG3;
wire[2-1:0] DEBUG_select_S4BEG0;
wire[2-1:0] DEBUG_select_S4BEG1;
wire[2-1:0] DEBUG_select_S4BEG2;
wire[2-1:0] DEBUG_select_S4BEG3;
wire[3-1:0] DEBUG_select_SS4BEG0;
wire[3-1:0] DEBUG_select_SS4BEG1;
wire[3-1:0] DEBUG_select_SS4BEG2;
wire[3-1:0] DEBUG_select_SS4BEG3;
wire[2-1:0] DEBUG_select_W1BEG0;
wire[2-1:0] DEBUG_select_W1BEG1;
wire[2-1:0] DEBUG_select_W1BEG2;
wire[2-1:0] DEBUG_select_W1BEG3;
wire[3-1:0] DEBUG_select_WW4BEG0;
wire[3-1:0] DEBUG_select_WW4BEG1;
wire[3-1:0] DEBUG_select_WW4BEG2;
wire[3-1:0] DEBUG_select_WW4BEG3;
wire[4-1:0] DEBUG_select_W6BEG0;
wire[4-1:0] DEBUG_select_W6BEG1;
wire[2-1:0] DEBUG_select_J2MID_ABa_BEG0;
wire[2-1:0] DEBUG_select_J2MID_ABa_BEG1;
wire[2-1:0] DEBUG_select_J2MID_ABa_BEG2;
wire[2-1:0] DEBUG_select_J2MID_ABa_BEG3;
wire[2-1:0] DEBUG_select_J2MID_CDa_BEG0;
wire[2-1:0] DEBUG_select_J2MID_CDa_BEG1;
wire[2-1:0] DEBUG_select_J2MID_CDa_BEG2;
wire[2-1:0] DEBUG_select_J2MID_CDa_BEG3;
wire[2-1:0] DEBUG_select_J2MID_EFa_BEG0;
wire[2-1:0] DEBUG_select_J2MID_EFa_BEG1;
wire[2-1:0] DEBUG_select_J2MID_EFa_BEG2;
wire[2-1:0] DEBUG_select_J2MID_EFa_BEG3;
wire[2-1:0] DEBUG_select_J2MID_GHa_BEG0;
wire[2-1:0] DEBUG_select_J2MID_GHa_BEG1;
wire[2-1:0] DEBUG_select_J2MID_GHa_BEG2;
wire[2-1:0] DEBUG_select_J2MID_GHa_BEG3;
wire[2-1:0] DEBUG_select_J2MID_ABb_BEG0;
wire[2-1:0] DEBUG_select_J2MID_ABb_BEG1;
wire[2-1:0] DEBUG_select_J2MID_ABb_BEG2;
wire[2-1:0] DEBUG_select_J2MID_ABb_BEG3;
wire[2-1:0] DEBUG_select_J2MID_CDb_BEG0;
wire[2-1:0] DEBUG_select_J2MID_CDb_BEG1;
wire[2-1:0] DEBUG_select_J2MID_CDb_BEG2;
wire[2-1:0] DEBUG_select_J2MID_CDb_BEG3;
wire[2-1:0] DEBUG_select_J2MID_EFb_BEG0;
wire[2-1:0] DEBUG_select_J2MID_EFb_BEG1;
wire[2-1:0] DEBUG_select_J2MID_EFb_BEG2;
wire[2-1:0] DEBUG_select_J2MID_EFb_BEG3;
wire[2-1:0] DEBUG_select_J2MID_GHb_BEG0;
wire[2-1:0] DEBUG_select_J2MID_GHb_BEG1;
wire[2-1:0] DEBUG_select_J2MID_GHb_BEG2;
wire[2-1:0] DEBUG_select_J2MID_GHb_BEG3;
wire[2-1:0] DEBUG_select_J2END_AB_BEG0;
wire[2-1:0] DEBUG_select_J2END_AB_BEG1;
wire[2-1:0] DEBUG_select_J2END_AB_BEG2;
wire[2-1:0] DEBUG_select_J2END_AB_BEG3;
wire[2-1:0] DEBUG_select_J2END_CD_BEG0;
wire[2-1:0] DEBUG_select_J2END_CD_BEG1;
wire[2-1:0] DEBUG_select_J2END_CD_BEG2;
wire[2-1:0] DEBUG_select_J2END_CD_BEG3;
wire[2-1:0] DEBUG_select_J2END_EF_BEG0;
wire[2-1:0] DEBUG_select_J2END_EF_BEG1;
wire[2-1:0] DEBUG_select_J2END_EF_BEG2;
wire[2-1:0] DEBUG_select_J2END_EF_BEG3;
wire[2-1:0] DEBUG_select_J2END_GH_BEG0;
wire[2-1:0] DEBUG_select_J2END_GH_BEG1;
wire[2-1:0] DEBUG_select_J2END_GH_BEG2;
wire[2-1:0] DEBUG_select_J2END_GH_BEG3;
wire[4-1:0] DEBUG_select_JN2BEG0;
wire[4-1:0] DEBUG_select_JN2BEG1;
wire[4-1:0] DEBUG_select_JN2BEG2;
wire[4-1:0] DEBUG_select_JN2BEG3;
wire[4-1:0] DEBUG_select_JN2BEG4;
wire[4-1:0] DEBUG_select_JN2BEG5;
wire[4-1:0] DEBUG_select_JN2BEG6;
wire[4-1:0] DEBUG_select_JN2BEG7;
wire[4-1:0] DEBUG_select_JE2BEG0;
wire[4-1:0] DEBUG_select_JE2BEG1;
wire[4-1:0] DEBUG_select_JE2BEG2;
wire[4-1:0] DEBUG_select_JE2BEG3;
wire[4-1:0] DEBUG_select_JE2BEG4;
wire[4-1:0] DEBUG_select_JE2BEG5;
wire[4-1:0] DEBUG_select_JE2BEG6;
wire[4-1:0] DEBUG_select_JE2BEG7;
wire[4-1:0] DEBUG_select_JS2BEG0;
wire[4-1:0] DEBUG_select_JS2BEG1;
wire[4-1:0] DEBUG_select_JS2BEG2;
wire[4-1:0] DEBUG_select_JS2BEG3;
wire[4-1:0] DEBUG_select_JS2BEG4;
wire[4-1:0] DEBUG_select_JS2BEG5;
wire[4-1:0] DEBUG_select_JS2BEG6;
wire[4-1:0] DEBUG_select_JS2BEG7;
wire[4-1:0] DEBUG_select_JW2BEG0;
wire[4-1:0] DEBUG_select_JW2BEG1;
wire[4-1:0] DEBUG_select_JW2BEG2;
wire[4-1:0] DEBUG_select_JW2BEG3;
wire[4-1:0] DEBUG_select_JW2BEG4;
wire[4-1:0] DEBUG_select_JW2BEG5;
wire[4-1:0] DEBUG_select_JW2BEG6;
wire[4-1:0] DEBUG_select_JW2BEG7;
wire[2-1:0] DEBUG_select_J_l_AB_BEG0;
wire[2-1:0] DEBUG_select_J_l_AB_BEG1;
wire[2-1:0] DEBUG_select_J_l_AB_BEG2;
wire[2-1:0] DEBUG_select_J_l_AB_BEG3;
wire[2-1:0] DEBUG_select_J_l_CD_BEG0;
wire[2-1:0] DEBUG_select_J_l_CD_BEG1;
wire[2-1:0] DEBUG_select_J_l_CD_BEG2;
wire[2-1:0] DEBUG_select_J_l_CD_BEG3;
wire[2-1:0] DEBUG_select_J_l_EF_BEG0;
wire[2-1:0] DEBUG_select_J_l_EF_BEG1;
wire[2-1:0] DEBUG_select_J_l_EF_BEG2;
wire[2-1:0] DEBUG_select_J_l_EF_BEG3;
wire[2-1:0] DEBUG_select_J_l_GH_BEG0;
wire[2-1:0] DEBUG_select_J_l_GH_BEG1;
wire[2-1:0] DEBUG_select_J_l_GH_BEG2;
wire[2-1:0] DEBUG_select_J_l_GH_BEG3;
 //The configuration bits (if any) are just a long shift register
 //This shift register is padded to an even number of flops/latches
 //switch matrix multiplexer i_2to60 MUX-4
assign i_2to60_input = {J_l_AB_END0,J2END_AB_END0,J2MID_ABb_END0,J2MID_ABa_END0};
cus_mux41_buf inst_cus_mux41_buf_i_2to60 (
    .A0(i_2to60_input[0]),
    .A1(i_2to60_input[1]),
    .A2(i_2to60_input[2]),
    .A3(i_2to60_input[3]),
    .S0(ConfigBits[0+0]),
    .S0N(ConfigBits_N[0+0]),
    .S1(ConfigBits[0+1]),
    .S1N(ConfigBits_N[0+1]),
    .X(i_2to60)
);

 //switch matrix multiplexer i_2to61 MUX-4
assign i_2to61_input = {J_l_AB_END1,J2END_AB_END1,J2MID_ABb_END1,J2MID_ABa_END1};
cus_mux41_buf inst_cus_mux41_buf_i_2to61 (
    .A0(i_2to61_input[0]),
    .A1(i_2to61_input[1]),
    .A2(i_2to61_input[2]),
    .A3(i_2to61_input[3]),
    .S0(ConfigBits[2+0]),
    .S0N(ConfigBits_N[2+0]),
    .S1(ConfigBits[2+1]),
    .S1N(ConfigBits_N[2+1]),
    .X(i_2to61)
);

 //switch matrix multiplexer i_2to62 MUX-4
assign i_2to62_input = {J_l_CD_END2,J2END_CD_END2,J2MID_CDb_END2,J2MID_CDa_END2};
cus_mux41_buf inst_cus_mux41_buf_i_2to62 (
    .A0(i_2to62_input[0]),
    .A1(i_2to62_input[1]),
    .A2(i_2to62_input[2]),
    .A3(i_2to62_input[3]),
    .S0(ConfigBits[4+0]),
    .S0N(ConfigBits_N[4+0]),
    .S1(ConfigBits[4+1]),
    .S1N(ConfigBits_N[4+1]),
    .X(i_2to62)
);

 //switch matrix multiplexer i_2to63 MUX-4
assign i_2to63_input = {J_l_CD_END3,J2END_CD_END3,J2MID_CDb_END3,J2MID_CDa_END3};
cus_mux41_buf inst_cus_mux41_buf_i_2to63 (
    .A0(i_2to63_input[0]),
    .A1(i_2to63_input[1]),
    .A2(i_2to63_input[2]),
    .A3(i_2to63_input[3]),
    .S0(ConfigBits[6+0]),
    .S0N(ConfigBits_N[6+0]),
    .S1(ConfigBits[6+1]),
    .S1N(ConfigBits_N[6+1]),
    .X(i_2to63)
);

 //switch matrix multiplexer i_2to64 MUX-4
assign i_2to64_input = {J_l_EF_END0,J2END_EF_END0,J2MID_EFb_END0,J2MID_EFa_END0};
cus_mux41_buf inst_cus_mux41_buf_i_2to64 (
    .A0(i_2to64_input[0]),
    .A1(i_2to64_input[1]),
    .A2(i_2to64_input[2]),
    .A3(i_2to64_input[3]),
    .S0(ConfigBits[8+0]),
    .S0N(ConfigBits_N[8+0]),
    .S1(ConfigBits[8+1]),
    .S1N(ConfigBits_N[8+1]),
    .X(i_2to64)
);

 //switch matrix multiplexer i_2to65 MUX-4
assign i_2to65_input = {J_l_EF_END0,J2END_EF_END0,J2MID_EFb_END0,J2MID_EFa_END0};
cus_mux41_buf inst_cus_mux41_buf_i_2to65 (
    .A0(i_2to65_input[0]),
    .A1(i_2to65_input[1]),
    .A2(i_2to65_input[2]),
    .A3(i_2to65_input[3]),
    .S0(ConfigBits[10+0]),
    .S0N(ConfigBits_N[10+0]),
    .S1(ConfigBits[10+1]),
    .S1N(ConfigBits_N[10+1]),
    .X(i_2to65)
);

 //switch matrix multiplexer i_2to66 MUX-4
assign i_2to66_input = {J_l_GH_END0,J2END_GH_END0,J2MID_GHb_END0,J2MID_GHa_END0};
cus_mux41_buf inst_cus_mux41_buf_i_2to66 (
    .A0(i_2to66_input[0]),
    .A1(i_2to66_input[1]),
    .A2(i_2to66_input[2]),
    .A3(i_2to66_input[3]),
    .S0(ConfigBits[12+0]),
    .S0N(ConfigBits_N[12+0]),
    .S1(ConfigBits[12+1]),
    .S1N(ConfigBits_N[12+1]),
    .X(i_2to66)
);

 //switch matrix multiplexer i_2to67 MUX-4
assign i_2to67_input = {J_l_GH_END0,J2END_GH_END0,J2MID_GHb_END0,J2MID_GHa_END0};
cus_mux41_buf inst_cus_mux41_buf_i_2to67 (
    .A0(i_2to67_input[0]),
    .A1(i_2to67_input[1]),
    .A2(i_2to67_input[2]),
    .A3(i_2to67_input[3]),
    .S0(ConfigBits[14+0]),
    .S0N(ConfigBits_N[14+0]),
    .S1(ConfigBits[14+1]),
    .S1N(ConfigBits_N[14+1]),
    .X(i_2to67)
);

 //switch matrix multiplexer i_2to68 MUX-0
 //WARNING unused multiplexer MUX-i_2to68
 //switch matrix multiplexer i_2to69 MUX-0
 //WARNING unused multiplexer MUX-i_2to69
 //switch matrix multiplexer i_2to610 MUX-0
 //WARNING unused multiplexer MUX-i_2to610
 //switch matrix multiplexer i_2to611 MUX-0
 //WARNING unused multiplexer MUX-i_2to611
 //switch matrix multiplexer i_2to612 MUX-0
 //WARNING unused multiplexer MUX-i_2to612
 //switch matrix multiplexer i_2to613 MUX-0
 //WARNING unused multiplexer MUX-i_2to613
 //switch matrix multiplexer i_2to614 MUX-0
 //WARNING unused multiplexer MUX-i_2to614
 //switch matrix multiplexer i_2to615 MUX-0
 //WARNING unused multiplexer MUX-i_2to615
 //switch matrix multiplexer i_2to616 MUX-0
 //WARNING unused multiplexer MUX-i_2to616
 //switch matrix multiplexer i_2to617 MUX-0
 //WARNING unused multiplexer MUX-i_2to617
 //switch matrix multiplexer i_2to618 MUX-0
 //WARNING unused multiplexer MUX-i_2to618
 //switch matrix multiplexer i_2to619 MUX-0
 //WARNING unused multiplexer MUX-i_2to619
 //switch matrix multiplexer i_2to620 MUX-0
 //WARNING unused multiplexer MUX-i_2to620
 //switch matrix multiplexer i_2to621 MUX-0
 //WARNING unused multiplexer MUX-i_2to621
 //switch matrix multiplexer i_2to622 MUX-0
 //WARNING unused multiplexer MUX-i_2to622
 //switch matrix multiplexer i_2to623 MUX-0
 //WARNING unused multiplexer MUX-i_2to623
 //switch matrix multiplexer i_2to624 MUX-0
 //WARNING unused multiplexer MUX-i_2to624
 //switch matrix multiplexer i_2to625 MUX-0
 //WARNING unused multiplexer MUX-i_2to625
 //switch matrix multiplexer i_2to626 MUX-0
 //WARNING unused multiplexer MUX-i_2to626
 //switch matrix multiplexer i_2to627 MUX-0
 //WARNING unused multiplexer MUX-i_2to627
 //switch matrix multiplexer i_2to628 MUX-0
 //WARNING unused multiplexer MUX-i_2to628
 //switch matrix multiplexer i_2to629 MUX-0
 //WARNING unused multiplexer MUX-i_2to629
 //switch matrix multiplexer i_2to630 MUX-0
 //WARNING unused multiplexer MUX-i_2to630
 //switch matrix multiplexer i_2to631 MUX-0
 //WARNING unused multiplexer MUX-i_2to631
 //switch matrix multiplexer N1BEG0 MUX-4
assign N1BEG0_input = {J_l_CD_END1,JW2END3,J2MID_CDb_END3,o_6to22};
cus_mux41_buf inst_cus_mux41_buf_N1BEG0 (
    .A0(N1BEG0_input[0]),
    .A1(N1BEG0_input[1]),
    .A2(N1BEG0_input[2]),
    .A3(N1BEG0_input[3]),
    .S0(ConfigBits[16+0]),
    .S0N(ConfigBits_N[16+0]),
    .S1(ConfigBits[16+1]),
    .S1N(ConfigBits_N[16+1]),
    .X(N1BEG0)
);

 //switch matrix multiplexer N1BEG1 MUX-4
assign N1BEG1_input = {J_l_EF_END2,JW2END0,J2MID_EFb_END0,o_6to23};
cus_mux41_buf inst_cus_mux41_buf_N1BEG1 (
    .A0(N1BEG1_input[0]),
    .A1(N1BEG1_input[1]),
    .A2(N1BEG1_input[2]),
    .A3(N1BEG1_input[3]),
    .S0(ConfigBits[18+0]),
    .S0N(ConfigBits_N[18+0]),
    .S1(ConfigBits[18+1]),
    .S1N(ConfigBits_N[18+1]),
    .X(N1BEG1)
);

 //switch matrix multiplexer N1BEG2 MUX-4
assign N1BEG2_input = {J_l_GH_END3,JW2END1,J2MID_GHb_END1,o_6to24};
cus_mux41_buf inst_cus_mux41_buf_N1BEG2 (
    .A0(N1BEG2_input[0]),
    .A1(N1BEG2_input[1]),
    .A2(N1BEG2_input[2]),
    .A3(N1BEG2_input[3]),
    .S0(ConfigBits[20+0]),
    .S0N(ConfigBits_N[20+0]),
    .S1(ConfigBits[20+1]),
    .S1N(ConfigBits_N[20+1]),
    .X(N1BEG2)
);

 //switch matrix multiplexer N1BEG3 MUX-4
assign N1BEG3_input = {J_l_AB_END0,JW2END2,J2MID_ABb_END2,o_6to25};
cus_mux41_buf inst_cus_mux41_buf_N1BEG3 (
    .A0(N1BEG3_input[0]),
    .A1(N1BEG3_input[1]),
    .A2(N1BEG3_input[2]),
    .A3(N1BEG3_input[3]),
    .S0(ConfigBits[22+0]),
    .S0N(ConfigBits_N[22+0]),
    .S1(ConfigBits[22+1]),
    .S1N(ConfigBits_N[22+1]),
    .X(N1BEG3)
);

 //switch matrix multiplexer N2BEG0 MUX-1
assign N2BEG0 = JN2END0;

 //switch matrix multiplexer N2BEG1 MUX-1
assign N2BEG1 = JN2END1;

 //switch matrix multiplexer N2BEG2 MUX-1
assign N2BEG2 = JN2END2;

 //switch matrix multiplexer N2BEG3 MUX-1
assign N2BEG3 = JN2END3;

 //switch matrix multiplexer N2BEG4 MUX-1
assign N2BEG4 = JN2END4;

 //switch matrix multiplexer N2BEG5 MUX-1
assign N2BEG5 = JN2END5;

 //switch matrix multiplexer N2BEG6 MUX-1
assign N2BEG6 = JN2END6;

 //switch matrix multiplexer N2BEG7 MUX-1
assign N2BEG7 = JN2END7;

 //switch matrix multiplexer N2BEGb0 MUX-1
assign N2BEGb0 = N2MID0;

 //switch matrix multiplexer N2BEGb1 MUX-1
assign N2BEGb1 = N2MID1;

 //switch matrix multiplexer N2BEGb2 MUX-1
assign N2BEGb2 = N2MID2;

 //switch matrix multiplexer N2BEGb3 MUX-1
assign N2BEGb3 = N2MID3;

 //switch matrix multiplexer N2BEGb4 MUX-1
assign N2BEGb4 = N2MID4;

 //switch matrix multiplexer N2BEGb5 MUX-1
assign N2BEGb5 = N2MID5;

 //switch matrix multiplexer N2BEGb6 MUX-1
assign N2BEGb6 = N2MID6;

 //switch matrix multiplexer N2BEGb7 MUX-1
assign N2BEGb7 = N2MID7;

 //switch matrix multiplexer N4BEG0 MUX-4
assign N4BEG0_input = {E6END1,N4END1,N2END2,o_6to24};
cus_mux41_buf inst_cus_mux41_buf_N4BEG0 (
    .A0(N4BEG0_input[0]),
    .A1(N4BEG0_input[1]),
    .A2(N4BEG0_input[2]),
    .A3(N4BEG0_input[3]),
    .S0(ConfigBits[24+0]),
    .S0N(ConfigBits_N[24+0]),
    .S1(ConfigBits[24+1]),
    .S1N(ConfigBits_N[24+1]),
    .X(N4BEG0)
);

 //switch matrix multiplexer N4BEG1 MUX-4
assign N4BEG1_input = {E6END0,N4END2,N2END3,o_6to25};
cus_mux41_buf inst_cus_mux41_buf_N4BEG1 (
    .A0(N4BEG1_input[0]),
    .A1(N4BEG1_input[1]),
    .A2(N4BEG1_input[2]),
    .A3(N4BEG1_input[3]),
    .S0(ConfigBits[26+0]),
    .S0N(ConfigBits_N[26+0]),
    .S1(ConfigBits[26+1]),
    .S1N(ConfigBits_N[26+1]),
    .X(N4BEG1)
);

 //switch matrix multiplexer N4BEG2 MUX-4
assign N4BEG2_input = {W6END1,N4END3,N2END0,o_6to26};
cus_mux41_buf inst_cus_mux41_buf_N4BEG2 (
    .A0(N4BEG2_input[0]),
    .A1(N4BEG2_input[1]),
    .A2(N4BEG2_input[2]),
    .A3(N4BEG2_input[3]),
    .S0(ConfigBits[28+0]),
    .S0N(ConfigBits_N[28+0]),
    .S1(ConfigBits[28+1]),
    .S1N(ConfigBits_N[28+1]),
    .X(N4BEG2)
);

 //switch matrix multiplexer N4BEG3 MUX-4
assign N4BEG3_input = {W6END0,N4END0,N2END1,o_6to27};
cus_mux41_buf inst_cus_mux41_buf_N4BEG3 (
    .A0(N4BEG3_input[0]),
    .A1(N4BEG3_input[1]),
    .A2(N4BEG3_input[2]),
    .A3(N4BEG3_input[3]),
    .S0(ConfigBits[30+0]),
    .S0N(ConfigBits_N[30+0]),
    .S1(ConfigBits[30+1]),
    .S1N(ConfigBits_N[30+1]),
    .X(N4BEG3)
);

 //switch matrix multiplexer NN4BEG0 MUX-8
assign NN4BEG0_input = {J2END_GH_END1,J2MID_CDb_END1,J2MID_ABb_END1,W1END2,E1END2,N1END2,o_6to26,o_6to25};
cus_mux81_buf inst_cus_mux81_buf_NN4BEG0 (
    .A0(NN4BEG0_input[0]),
    .A1(NN4BEG0_input[1]),
    .A2(NN4BEG0_input[2]),
    .A3(NN4BEG0_input[3]),
    .A4(NN4BEG0_input[4]),
    .A5(NN4BEG0_input[5]),
    .A6(NN4BEG0_input[6]),
    .A7(NN4BEG0_input[7]),
    .S0(ConfigBits[32+0]),
    .S0N(ConfigBits_N[32+0]),
    .S1(ConfigBits[32+1]),
    .S1N(ConfigBits_N[32+1]),
    .S2(ConfigBits[32+2]),
    .S2N(ConfigBits_N[32+2]),
    .X(NN4BEG0)
);

 //switch matrix multiplexer NN4BEG1 MUX-8
assign NN4BEG1_input = {J2END_EF_END1,J2MID_CDa_END2,J2MID_ABa_END2,W1END3,E1END3,N1END3,o_6to27,o_6to20};
cus_mux81_buf inst_cus_mux81_buf_NN4BEG1 (
    .A0(NN4BEG1_input[0]),
    .A1(NN4BEG1_input[1]),
    .A2(NN4BEG1_input[2]),
    .A3(NN4BEG1_input[3]),
    .A4(NN4BEG1_input[4]),
    .A5(NN4BEG1_input[5]),
    .A6(NN4BEG1_input[6]),
    .A7(NN4BEG1_input[7]),
    .S0(ConfigBits[35+0]),
    .S0N(ConfigBits_N[35+0]),
    .S1(ConfigBits[35+1]),
    .S1N(ConfigBits_N[35+1]),
    .S2(ConfigBits[35+2]),
    .S2N(ConfigBits_N[35+2]),
    .X(NN4BEG1)
);

 //switch matrix multiplexer NN4BEG2 MUX-8
assign NN4BEG2_input = {J2END_CD_END1,J2MID_GHb_END1,J2MID_EFb_END1,W1END0,E1END0,N1END0,o_6to22,o_6to21};
cus_mux81_buf inst_cus_mux81_buf_NN4BEG2 (
    .A0(NN4BEG2_input[0]),
    .A1(NN4BEG2_input[1]),
    .A2(NN4BEG2_input[2]),
    .A3(NN4BEG2_input[3]),
    .A4(NN4BEG2_input[4]),
    .A5(NN4BEG2_input[5]),
    .A6(NN4BEG2_input[6]),
    .A7(NN4BEG2_input[7]),
    .S0(ConfigBits[38+0]),
    .S0N(ConfigBits_N[38+0]),
    .S1(ConfigBits[38+1]),
    .S1N(ConfigBits_N[38+1]),
    .S2(ConfigBits[38+2]),
    .S2N(ConfigBits_N[38+2]),
    .X(NN4BEG2)
);

 //switch matrix multiplexer NN4BEG3 MUX-8
assign NN4BEG3_input = {J2END_AB_END1,J2MID_GHa_END2,J2MID_EFa_END2,W1END1,E1END1,N1END1,o_6to24,o_6to23};
cus_mux81_buf inst_cus_mux81_buf_NN4BEG3 (
    .A0(NN4BEG3_input[0]),
    .A1(NN4BEG3_input[1]),
    .A2(NN4BEG3_input[2]),
    .A3(NN4BEG3_input[3]),
    .A4(NN4BEG3_input[4]),
    .A5(NN4BEG3_input[5]),
    .A6(NN4BEG3_input[6]),
    .A7(NN4BEG3_input[7]),
    .S0(ConfigBits[41+0]),
    .S0N(ConfigBits_N[41+0]),
    .S1(ConfigBits[41+1]),
    .S1N(ConfigBits_N[41+1]),
    .S2(ConfigBits[41+2]),
    .S2N(ConfigBits_N[41+2]),
    .X(NN4BEG3)
);

 //switch matrix multiplexer E1BEG0 MUX-4
assign E1BEG0_input = {J_l_CD_END1,JN2END3,J2MID_CDb_END3,o_6to23};
cus_mux41_buf inst_cus_mux41_buf_E1BEG0 (
    .A0(E1BEG0_input[0]),
    .A1(E1BEG0_input[1]),
    .A2(E1BEG0_input[2]),
    .A3(E1BEG0_input[3]),
    .S0(ConfigBits[44+0]),
    .S0N(ConfigBits_N[44+0]),
    .S1(ConfigBits[44+1]),
    .S1N(ConfigBits_N[44+1]),
    .X(E1BEG0)
);

 //switch matrix multiplexer E1BEG1 MUX-4
assign E1BEG1_input = {J_l_EF_END2,JN2END0,J2MID_EFb_END0,o_6to24};
cus_mux41_buf inst_cus_mux41_buf_E1BEG1 (
    .A0(E1BEG1_input[0]),
    .A1(E1BEG1_input[1]),
    .A2(E1BEG1_input[2]),
    .A3(E1BEG1_input[3]),
    .S0(ConfigBits[46+0]),
    .S0N(ConfigBits_N[46+0]),
    .S1(ConfigBits[46+1]),
    .S1N(ConfigBits_N[46+1]),
    .X(E1BEG1)
);

 //switch matrix multiplexer E1BEG2 MUX-4
assign E1BEG2_input = {J_l_GH_END3,JN2END1,J2MID_GHb_END1,o_6to25};
cus_mux41_buf inst_cus_mux41_buf_E1BEG2 (
    .A0(E1BEG2_input[0]),
    .A1(E1BEG2_input[1]),
    .A2(E1BEG2_input[2]),
    .A3(E1BEG2_input[3]),
    .S0(ConfigBits[48+0]),
    .S0N(ConfigBits_N[48+0]),
    .S1(ConfigBits[48+1]),
    .S1N(ConfigBits_N[48+1]),
    .X(E1BEG2)
);

 //switch matrix multiplexer E1BEG3 MUX-4
assign E1BEG3_input = {J_l_AB_END0,JN2END2,J2MID_ABb_END2,o_6to26};
cus_mux41_buf inst_cus_mux41_buf_E1BEG3 (
    .A0(E1BEG3_input[0]),
    .A1(E1BEG3_input[1]),
    .A2(E1BEG3_input[2]),
    .A3(E1BEG3_input[3]),
    .S0(ConfigBits[50+0]),
    .S0N(ConfigBits_N[50+0]),
    .S1(ConfigBits[50+1]),
    .S1N(ConfigBits_N[50+1]),
    .X(E1BEG3)
);

 //switch matrix multiplexer E2BEG0 MUX-1
assign E2BEG0 = JE2END0;

 //switch matrix multiplexer E2BEG1 MUX-1
assign E2BEG1 = JE2END1;

 //switch matrix multiplexer E2BEG2 MUX-1
assign E2BEG2 = JE2END2;

 //switch matrix multiplexer E2BEG3 MUX-1
assign E2BEG3 = JE2END3;

 //switch matrix multiplexer E2BEG4 MUX-1
assign E2BEG4 = JE2END4;

 //switch matrix multiplexer E2BEG5 MUX-1
assign E2BEG5 = JE2END5;

 //switch matrix multiplexer E2BEG6 MUX-1
assign E2BEG6 = JE2END6;

 //switch matrix multiplexer E2BEG7 MUX-1
assign E2BEG7 = JE2END7;

 //switch matrix multiplexer E2BEGb0 MUX-1
assign E2BEGb0 = E2MID0;

 //switch matrix multiplexer E2BEGb1 MUX-1
assign E2BEGb1 = E2MID1;

 //switch matrix multiplexer E2BEGb2 MUX-1
assign E2BEGb2 = E2MID2;

 //switch matrix multiplexer E2BEGb3 MUX-1
assign E2BEGb3 = E2MID3;

 //switch matrix multiplexer E2BEGb4 MUX-1
assign E2BEGb4 = E2MID4;

 //switch matrix multiplexer E2BEGb5 MUX-1
assign E2BEGb5 = E2MID5;

 //switch matrix multiplexer E2BEGb6 MUX-1
assign E2BEGb6 = E2MID6;

 //switch matrix multiplexer E2BEGb7 MUX-1
assign E2BEGb7 = E2MID7;

 //switch matrix multiplexer EE4BEG0 MUX-8
assign EE4BEG0_input = {J2END_GH_END0,J2MID_CDb_END1,J2MID_ABb_END1,S1END2,E1END2,N1END2,o_6to26,o_6to25};
cus_mux81_buf inst_cus_mux81_buf_EE4BEG0 (
    .A0(EE4BEG0_input[0]),
    .A1(EE4BEG0_input[1]),
    .A2(EE4BEG0_input[2]),
    .A3(EE4BEG0_input[3]),
    .A4(EE4BEG0_input[4]),
    .A5(EE4BEG0_input[5]),
    .A6(EE4BEG0_input[6]),
    .A7(EE4BEG0_input[7]),
    .S0(ConfigBits[52+0]),
    .S0N(ConfigBits_N[52+0]),
    .S1(ConfigBits[52+1]),
    .S1N(ConfigBits_N[52+1]),
    .S2(ConfigBits[52+2]),
    .S2N(ConfigBits_N[52+2]),
    .X(EE4BEG0)
);

 //switch matrix multiplexer EE4BEG1 MUX-8
assign EE4BEG1_input = {J2END_EF_END0,J2MID_CDa_END2,J2MID_ABa_END2,S1END3,E1END3,N1END3,o_6to27,o_6to20};
cus_mux81_buf inst_cus_mux81_buf_EE4BEG1 (
    .A0(EE4BEG1_input[0]),
    .A1(EE4BEG1_input[1]),
    .A2(EE4BEG1_input[2]),
    .A3(EE4BEG1_input[3]),
    .A4(EE4BEG1_input[4]),
    .A5(EE4BEG1_input[5]),
    .A6(EE4BEG1_input[6]),
    .A7(EE4BEG1_input[7]),
    .S0(ConfigBits[55+0]),
    .S0N(ConfigBits_N[55+0]),
    .S1(ConfigBits[55+1]),
    .S1N(ConfigBits_N[55+1]),
    .S2(ConfigBits[55+2]),
    .S2N(ConfigBits_N[55+2]),
    .X(EE4BEG1)
);

 //switch matrix multiplexer EE4BEG2 MUX-8
assign EE4BEG2_input = {J2END_CD_END0,J2MID_GHb_END1,J2MID_EFb_END1,S1END0,E1END0,N1END0,o_6to22,o_6to21};
cus_mux81_buf inst_cus_mux81_buf_EE4BEG2 (
    .A0(EE4BEG2_input[0]),
    .A1(EE4BEG2_input[1]),
    .A2(EE4BEG2_input[2]),
    .A3(EE4BEG2_input[3]),
    .A4(EE4BEG2_input[4]),
    .A5(EE4BEG2_input[5]),
    .A6(EE4BEG2_input[6]),
    .A7(EE4BEG2_input[7]),
    .S0(ConfigBits[58+0]),
    .S0N(ConfigBits_N[58+0]),
    .S1(ConfigBits[58+1]),
    .S1N(ConfigBits_N[58+1]),
    .S2(ConfigBits[58+2]),
    .S2N(ConfigBits_N[58+2]),
    .X(EE4BEG2)
);

 //switch matrix multiplexer EE4BEG3 MUX-8
assign EE4BEG3_input = {J2END_AB_END0,J2MID_GHa_END2,J2MID_EFa_END2,S1END1,E1END1,N1END1,o_6to24,o_6to23};
cus_mux81_buf inst_cus_mux81_buf_EE4BEG3 (
    .A0(EE4BEG3_input[0]),
    .A1(EE4BEG3_input[1]),
    .A2(EE4BEG3_input[2]),
    .A3(EE4BEG3_input[3]),
    .A4(EE4BEG3_input[4]),
    .A5(EE4BEG3_input[5]),
    .A6(EE4BEG3_input[6]),
    .A7(EE4BEG3_input[7]),
    .S0(ConfigBits[61+0]),
    .S0N(ConfigBits_N[61+0]),
    .S1(ConfigBits[61+1]),
    .S1N(ConfigBits_N[61+1]),
    .S2(ConfigBits[61+2]),
    .S2N(ConfigBits_N[61+2]),
    .X(EE4BEG3)
);

 //switch matrix multiplexer E6BEG0 MUX-16
assign E6BEG0_input = {J2MID_GHb_END1,J2MID_EFb_END1,J2MID_CDb_END1,J2MID_ABb_END1,W1END3,SS4END0,E1END3,NN4END0,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_E6BEG0 (
    .A0(E6BEG0_input[0]),
    .A1(E6BEG0_input[1]),
    .A2(E6BEG0_input[2]),
    .A3(E6BEG0_input[3]),
    .A4(E6BEG0_input[4]),
    .A5(E6BEG0_input[5]),
    .A6(E6BEG0_input[6]),
    .A7(E6BEG0_input[7]),
    .A8(E6BEG0_input[8]),
    .A9(E6BEG0_input[9]),
    .A10(E6BEG0_input[10]),
    .A11(E6BEG0_input[11]),
    .A12(E6BEG0_input[12]),
    .A13(E6BEG0_input[13]),
    .A14(E6BEG0_input[14]),
    .A15(E6BEG0_input[15]),
    .S0(ConfigBits[64+0]),
    .S0N(ConfigBits_N[64+0]),
    .S1(ConfigBits[64+1]),
    .S1N(ConfigBits_N[64+1]),
    .S2(ConfigBits[64+2]),
    .S2N(ConfigBits_N[64+2]),
    .S3(ConfigBits[64+3]),
    .S3N(ConfigBits_N[64+3]),
    .X(E6BEG0)
);

 //switch matrix multiplexer E6BEG1 MUX-16
assign E6BEG1_input = {J2MID_GHa_END2,J2MID_EFa_END2,J2MID_CDa_END2,J2MID_ABa_END2,W1END2,SS4END3,E1END2,NN4END3,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_E6BEG1 (
    .A0(E6BEG1_input[0]),
    .A1(E6BEG1_input[1]),
    .A2(E6BEG1_input[2]),
    .A3(E6BEG1_input[3]),
    .A4(E6BEG1_input[4]),
    .A5(E6BEG1_input[5]),
    .A6(E6BEG1_input[6]),
    .A7(E6BEG1_input[7]),
    .A8(E6BEG1_input[8]),
    .A9(E6BEG1_input[9]),
    .A10(E6BEG1_input[10]),
    .A11(E6BEG1_input[11]),
    .A12(E6BEG1_input[12]),
    .A13(E6BEG1_input[13]),
    .A14(E6BEG1_input[14]),
    .A15(E6BEG1_input[15]),
    .S0(ConfigBits[68+0]),
    .S0N(ConfigBits_N[68+0]),
    .S1(ConfigBits[68+1]),
    .S1N(ConfigBits_N[68+1]),
    .S2(ConfigBits[68+2]),
    .S2N(ConfigBits_N[68+2]),
    .S3(ConfigBits[68+3]),
    .S3N(ConfigBits_N[68+3]),
    .X(E6BEG1)
);

 //switch matrix multiplexer S1BEG0 MUX-4
assign S1BEG0_input = {J_l_CD_END1,JE2END3,J2MID_CDb_END3,o_6to24};
cus_mux41_buf inst_cus_mux41_buf_S1BEG0 (
    .A0(S1BEG0_input[0]),
    .A1(S1BEG0_input[1]),
    .A2(S1BEG0_input[2]),
    .A3(S1BEG0_input[3]),
    .S0(ConfigBits[72+0]),
    .S0N(ConfigBits_N[72+0]),
    .S1(ConfigBits[72+1]),
    .S1N(ConfigBits_N[72+1]),
    .X(S1BEG0)
);

 //switch matrix multiplexer S1BEG1 MUX-4
assign S1BEG1_input = {J_l_EF_END2,JE2END0,J2MID_EFb_END0,o_6to25};
cus_mux41_buf inst_cus_mux41_buf_S1BEG1 (
    .A0(S1BEG1_input[0]),
    .A1(S1BEG1_input[1]),
    .A2(S1BEG1_input[2]),
    .A3(S1BEG1_input[3]),
    .S0(ConfigBits[74+0]),
    .S0N(ConfigBits_N[74+0]),
    .S1(ConfigBits[74+1]),
    .S1N(ConfigBits_N[74+1]),
    .X(S1BEG1)
);

 //switch matrix multiplexer S1BEG2 MUX-4
assign S1BEG2_input = {J_l_GH_END3,JE2END1,J2MID_GHb_END1,o_6to26};
cus_mux41_buf inst_cus_mux41_buf_S1BEG2 (
    .A0(S1BEG2_input[0]),
    .A1(S1BEG2_input[1]),
    .A2(S1BEG2_input[2]),
    .A3(S1BEG2_input[3]),
    .S0(ConfigBits[76+0]),
    .S0N(ConfigBits_N[76+0]),
    .S1(ConfigBits[76+1]),
    .S1N(ConfigBits_N[76+1]),
    .X(S1BEG2)
);

 //switch matrix multiplexer S1BEG3 MUX-4
assign S1BEG3_input = {J_l_AB_END0,JE2END2,J2MID_ABb_END2,o_6to27};
cus_mux41_buf inst_cus_mux41_buf_S1BEG3 (
    .A0(S1BEG3_input[0]),
    .A1(S1BEG3_input[1]),
    .A2(S1BEG3_input[2]),
    .A3(S1BEG3_input[3]),
    .S0(ConfigBits[78+0]),
    .S0N(ConfigBits_N[78+0]),
    .S1(ConfigBits[78+1]),
    .S1N(ConfigBits_N[78+1]),
    .X(S1BEG3)
);

 //switch matrix multiplexer S2BEG0 MUX-1
assign S2BEG0 = JS2END0;

 //switch matrix multiplexer S2BEG1 MUX-1
assign S2BEG1 = JS2END1;

 //switch matrix multiplexer S2BEG2 MUX-1
assign S2BEG2 = JS2END2;

 //switch matrix multiplexer S2BEG3 MUX-1
assign S2BEG3 = JS2END3;

 //switch matrix multiplexer S2BEG4 MUX-1
assign S2BEG4 = JS2END4;

 //switch matrix multiplexer S2BEG5 MUX-1
assign S2BEG5 = JS2END5;

 //switch matrix multiplexer S2BEG6 MUX-1
assign S2BEG6 = JS2END6;

 //switch matrix multiplexer S2BEG7 MUX-1
assign S2BEG7 = JS2END7;

 //switch matrix multiplexer S2BEGb0 MUX-1
assign S2BEGb0 = S2MID0;

 //switch matrix multiplexer S2BEGb1 MUX-1
assign S2BEGb1 = S2MID1;

 //switch matrix multiplexer S2BEGb2 MUX-1
assign S2BEGb2 = S2MID2;

 //switch matrix multiplexer S2BEGb3 MUX-1
assign S2BEGb3 = S2MID3;

 //switch matrix multiplexer S2BEGb4 MUX-1
assign S2BEGb4 = S2MID4;

 //switch matrix multiplexer S2BEGb5 MUX-1
assign S2BEGb5 = S2MID5;

 //switch matrix multiplexer S2BEGb6 MUX-1
assign S2BEGb6 = S2MID6;

 //switch matrix multiplexer S2BEGb7 MUX-1
assign S2BEGb7 = S2MID7;

 //switch matrix multiplexer S4BEG0 MUX-4
assign S4BEG0_input = {S4END1,S2END2,E6END1,o_6to20};
cus_mux41_buf inst_cus_mux41_buf_S4BEG0 (
    .A0(S4BEG0_input[0]),
    .A1(S4BEG0_input[1]),
    .A2(S4BEG0_input[2]),
    .A3(S4BEG0_input[3]),
    .S0(ConfigBits[80+0]),
    .S0N(ConfigBits_N[80+0]),
    .S1(ConfigBits[80+1]),
    .S1N(ConfigBits_N[80+1]),
    .X(S4BEG0)
);

 //switch matrix multiplexer S4BEG1 MUX-4
assign S4BEG1_input = {S4END2,S2END3,E6END0,o_6to21};
cus_mux41_buf inst_cus_mux41_buf_S4BEG1 (
    .A0(S4BEG1_input[0]),
    .A1(S4BEG1_input[1]),
    .A2(S4BEG1_input[2]),
    .A3(S4BEG1_input[3]),
    .S0(ConfigBits[82+0]),
    .S0N(ConfigBits_N[82+0]),
    .S1(ConfigBits[82+1]),
    .S1N(ConfigBits_N[82+1]),
    .X(S4BEG1)
);

 //switch matrix multiplexer S4BEG2 MUX-4
assign S4BEG2_input = {W6END1,S4END3,S2END0,o_6to22};
cus_mux41_buf inst_cus_mux41_buf_S4BEG2 (
    .A0(S4BEG2_input[0]),
    .A1(S4BEG2_input[1]),
    .A2(S4BEG2_input[2]),
    .A3(S4BEG2_input[3]),
    .S0(ConfigBits[84+0]),
    .S0N(ConfigBits_N[84+0]),
    .S1(ConfigBits[84+1]),
    .S1N(ConfigBits_N[84+1]),
    .X(S4BEG2)
);

 //switch matrix multiplexer S4BEG3 MUX-4
assign S4BEG3_input = {W6END0,S4END0,S2END1,o_6to23};
cus_mux41_buf inst_cus_mux41_buf_S4BEG3 (
    .A0(S4BEG3_input[0]),
    .A1(S4BEG3_input[1]),
    .A2(S4BEG3_input[2]),
    .A3(S4BEG3_input[3]),
    .S0(ConfigBits[86+0]),
    .S0N(ConfigBits_N[86+0]),
    .S1(ConfigBits[86+1]),
    .S1N(ConfigBits_N[86+1]),
    .X(S4BEG3)
);

 //switch matrix multiplexer SS4BEG0 MUX-8
assign SS4BEG0_input = {J2END_GH_END3,J2MID_CDb_END1,J2MID_ABb_END1,W1END2,E1END2,N1END2,o_6to26,o_6to25};
cus_mux81_buf inst_cus_mux81_buf_SS4BEG0 (
    .A0(SS4BEG0_input[0]),
    .A1(SS4BEG0_input[1]),
    .A2(SS4BEG0_input[2]),
    .A3(SS4BEG0_input[3]),
    .A4(SS4BEG0_input[4]),
    .A5(SS4BEG0_input[5]),
    .A6(SS4BEG0_input[6]),
    .A7(SS4BEG0_input[7]),
    .S0(ConfigBits[88+0]),
    .S0N(ConfigBits_N[88+0]),
    .S1(ConfigBits[88+1]),
    .S1N(ConfigBits_N[88+1]),
    .S2(ConfigBits[88+2]),
    .S2N(ConfigBits_N[88+2]),
    .X(SS4BEG0)
);

 //switch matrix multiplexer SS4BEG1 MUX-8
assign SS4BEG1_input = {J2END_EF_END3,J2MID_CDa_END2,J2MID_ABa_END2,W1END3,E1END3,N1END3,o_6to27,o_6to20};
cus_mux81_buf inst_cus_mux81_buf_SS4BEG1 (
    .A0(SS4BEG1_input[0]),
    .A1(SS4BEG1_input[1]),
    .A2(SS4BEG1_input[2]),
    .A3(SS4BEG1_input[3]),
    .A4(SS4BEG1_input[4]),
    .A5(SS4BEG1_input[5]),
    .A6(SS4BEG1_input[6]),
    .A7(SS4BEG1_input[7]),
    .S0(ConfigBits[91+0]),
    .S0N(ConfigBits_N[91+0]),
    .S1(ConfigBits[91+1]),
    .S1N(ConfigBits_N[91+1]),
    .S2(ConfigBits[91+2]),
    .S2N(ConfigBits_N[91+2]),
    .X(SS4BEG1)
);

 //switch matrix multiplexer SS4BEG2 MUX-8
assign SS4BEG2_input = {J2END_CD_END3,J2MID_GHb_END1,J2MID_EFb_END1,W1END0,E1END0,N1END0,o_6to22,o_6to21};
cus_mux81_buf inst_cus_mux81_buf_SS4BEG2 (
    .A0(SS4BEG2_input[0]),
    .A1(SS4BEG2_input[1]),
    .A2(SS4BEG2_input[2]),
    .A3(SS4BEG2_input[3]),
    .A4(SS4BEG2_input[4]),
    .A5(SS4BEG2_input[5]),
    .A6(SS4BEG2_input[6]),
    .A7(SS4BEG2_input[7]),
    .S0(ConfigBits[94+0]),
    .S0N(ConfigBits_N[94+0]),
    .S1(ConfigBits[94+1]),
    .S1N(ConfigBits_N[94+1]),
    .S2(ConfigBits[94+2]),
    .S2N(ConfigBits_N[94+2]),
    .X(SS4BEG2)
);

 //switch matrix multiplexer SS4BEG3 MUX-8
assign SS4BEG3_input = {J2END_AB_END3,J2MID_GHa_END2,J2MID_EFa_END2,W1END1,E1END1,N1END1,o_6to24,o_6to23};
cus_mux81_buf inst_cus_mux81_buf_SS4BEG3 (
    .A0(SS4BEG3_input[0]),
    .A1(SS4BEG3_input[1]),
    .A2(SS4BEG3_input[2]),
    .A3(SS4BEG3_input[3]),
    .A4(SS4BEG3_input[4]),
    .A5(SS4BEG3_input[5]),
    .A6(SS4BEG3_input[6]),
    .A7(SS4BEG3_input[7]),
    .S0(ConfigBits[97+0]),
    .S0N(ConfigBits_N[97+0]),
    .S1(ConfigBits[97+1]),
    .S1N(ConfigBits_N[97+1]),
    .S2(ConfigBits[97+2]),
    .S2N(ConfigBits_N[97+2]),
    .X(SS4BEG3)
);

 //switch matrix multiplexer W1BEG0 MUX-4
assign W1BEG0_input = {J_l_CD_END1,JS2END3,J2MID_CDb_END3,o_6to25};
cus_mux41_buf inst_cus_mux41_buf_W1BEG0 (
    .A0(W1BEG0_input[0]),
    .A1(W1BEG0_input[1]),
    .A2(W1BEG0_input[2]),
    .A3(W1BEG0_input[3]),
    .S0(ConfigBits[100+0]),
    .S0N(ConfigBits_N[100+0]),
    .S1(ConfigBits[100+1]),
    .S1N(ConfigBits_N[100+1]),
    .X(W1BEG0)
);

 //switch matrix multiplexer W1BEG1 MUX-4
assign W1BEG1_input = {J_l_EF_END2,JS2END0,J2MID_EFb_END0,o_6to26};
cus_mux41_buf inst_cus_mux41_buf_W1BEG1 (
    .A0(W1BEG1_input[0]),
    .A1(W1BEG1_input[1]),
    .A2(W1BEG1_input[2]),
    .A3(W1BEG1_input[3]),
    .S0(ConfigBits[102+0]),
    .S0N(ConfigBits_N[102+0]),
    .S1(ConfigBits[102+1]),
    .S1N(ConfigBits_N[102+1]),
    .X(W1BEG1)
);

 //switch matrix multiplexer W1BEG2 MUX-4
assign W1BEG2_input = {J_l_GH_END3,JS2END1,J2MID_GHb_END1,o_6to27};
cus_mux41_buf inst_cus_mux41_buf_W1BEG2 (
    .A0(W1BEG2_input[0]),
    .A1(W1BEG2_input[1]),
    .A2(W1BEG2_input[2]),
    .A3(W1BEG2_input[3]),
    .S0(ConfigBits[104+0]),
    .S0N(ConfigBits_N[104+0]),
    .S1(ConfigBits[104+1]),
    .S1N(ConfigBits_N[104+1]),
    .X(W1BEG2)
);

 //switch matrix multiplexer W1BEG3 MUX-4
assign W1BEG3_input = {J_l_AB_END0,JS2END2,J2MID_ABb_END2,o_6to20};
cus_mux41_buf inst_cus_mux41_buf_W1BEG3 (
    .A0(W1BEG3_input[0]),
    .A1(W1BEG3_input[1]),
    .A2(W1BEG3_input[2]),
    .A3(W1BEG3_input[3]),
    .S0(ConfigBits[106+0]),
    .S0N(ConfigBits_N[106+0]),
    .S1(ConfigBits[106+1]),
    .S1N(ConfigBits_N[106+1]),
    .X(W1BEG3)
);

 //switch matrix multiplexer W2BEG0 MUX-1
assign W2BEG0 = JW2END0;

 //switch matrix multiplexer W2BEG1 MUX-1
assign W2BEG1 = JW2END1;

 //switch matrix multiplexer W2BEG2 MUX-1
assign W2BEG2 = JW2END2;

 //switch matrix multiplexer W2BEG3 MUX-1
assign W2BEG3 = JW2END3;

 //switch matrix multiplexer W2BEG4 MUX-1
assign W2BEG4 = JW2END4;

 //switch matrix multiplexer W2BEG5 MUX-1
assign W2BEG5 = JW2END5;

 //switch matrix multiplexer W2BEG6 MUX-1
assign W2BEG6 = JW2END6;

 //switch matrix multiplexer W2BEG7 MUX-1
assign W2BEG7 = JW2END7;

 //switch matrix multiplexer W2BEGb0 MUX-1
assign W2BEGb0 = W2MID0;

 //switch matrix multiplexer W2BEGb1 MUX-1
assign W2BEGb1 = W2MID1;

 //switch matrix multiplexer W2BEGb2 MUX-1
assign W2BEGb2 = W2MID2;

 //switch matrix multiplexer W2BEGb3 MUX-1
assign W2BEGb3 = W2MID3;

 //switch matrix multiplexer W2BEGb4 MUX-1
assign W2BEGb4 = W2MID4;

 //switch matrix multiplexer W2BEGb5 MUX-1
assign W2BEGb5 = W2MID5;

 //switch matrix multiplexer W2BEGb6 MUX-1
assign W2BEGb6 = W2MID6;

 //switch matrix multiplexer W2BEGb7 MUX-1
assign W2BEGb7 = W2MID7;

 //switch matrix multiplexer WW4BEG0 MUX-8
assign WW4BEG0_input = {J2END_GH_END2,J2MID_CDb_END1,J2MID_ABb_END1,W1END2,S1END2,N1END2,o_6to26,o_6to25};
cus_mux81_buf inst_cus_mux81_buf_WW4BEG0 (
    .A0(WW4BEG0_input[0]),
    .A1(WW4BEG0_input[1]),
    .A2(WW4BEG0_input[2]),
    .A3(WW4BEG0_input[3]),
    .A4(WW4BEG0_input[4]),
    .A5(WW4BEG0_input[5]),
    .A6(WW4BEG0_input[6]),
    .A7(WW4BEG0_input[7]),
    .S0(ConfigBits[108+0]),
    .S0N(ConfigBits_N[108+0]),
    .S1(ConfigBits[108+1]),
    .S1N(ConfigBits_N[108+1]),
    .S2(ConfigBits[108+2]),
    .S2N(ConfigBits_N[108+2]),
    .X(WW4BEG0)
);

 //switch matrix multiplexer WW4BEG1 MUX-8
assign WW4BEG1_input = {J2END_EF_END2,J2MID_CDa_END2,J2MID_ABa_END2,W1END3,S1END3,N1END3,o_6to27,o_6to20};
cus_mux81_buf inst_cus_mux81_buf_WW4BEG1 (
    .A0(WW4BEG1_input[0]),
    .A1(WW4BEG1_input[1]),
    .A2(WW4BEG1_input[2]),
    .A3(WW4BEG1_input[3]),
    .A4(WW4BEG1_input[4]),
    .A5(WW4BEG1_input[5]),
    .A6(WW4BEG1_input[6]),
    .A7(WW4BEG1_input[7]),
    .S0(ConfigBits[111+0]),
    .S0N(ConfigBits_N[111+0]),
    .S1(ConfigBits[111+1]),
    .S1N(ConfigBits_N[111+1]),
    .S2(ConfigBits[111+2]),
    .S2N(ConfigBits_N[111+2]),
    .X(WW4BEG1)
);

 //switch matrix multiplexer WW4BEG2 MUX-8
assign WW4BEG2_input = {J2END_CD_END2,J2MID_GHb_END1,J2MID_EFb_END1,W1END0,S1END0,N1END0,o_6to22,o_6to21};
cus_mux81_buf inst_cus_mux81_buf_WW4BEG2 (
    .A0(WW4BEG2_input[0]),
    .A1(WW4BEG2_input[1]),
    .A2(WW4BEG2_input[2]),
    .A3(WW4BEG2_input[3]),
    .A4(WW4BEG2_input[4]),
    .A5(WW4BEG2_input[5]),
    .A6(WW4BEG2_input[6]),
    .A7(WW4BEG2_input[7]),
    .S0(ConfigBits[114+0]),
    .S0N(ConfigBits_N[114+0]),
    .S1(ConfigBits[114+1]),
    .S1N(ConfigBits_N[114+1]),
    .S2(ConfigBits[114+2]),
    .S2N(ConfigBits_N[114+2]),
    .X(WW4BEG2)
);

 //switch matrix multiplexer WW4BEG3 MUX-8
assign WW4BEG3_input = {J2END_AB_END2,J2MID_GHa_END2,J2MID_EFa_END2,W1END1,S1END1,N1END1,o_6to24,o_6to23};
cus_mux81_buf inst_cus_mux81_buf_WW4BEG3 (
    .A0(WW4BEG3_input[0]),
    .A1(WW4BEG3_input[1]),
    .A2(WW4BEG3_input[2]),
    .A3(WW4BEG3_input[3]),
    .A4(WW4BEG3_input[4]),
    .A5(WW4BEG3_input[5]),
    .A6(WW4BEG3_input[6]),
    .A7(WW4BEG3_input[7]),
    .S0(ConfigBits[117+0]),
    .S0N(ConfigBits_N[117+0]),
    .S1(ConfigBits[117+1]),
    .S1N(ConfigBits_N[117+1]),
    .S2(ConfigBits[117+2]),
    .S2N(ConfigBits_N[117+2]),
    .X(WW4BEG3)
);

 //switch matrix multiplexer W6BEG0 MUX-16
assign W6BEG0_input = {J2MID_GHb_END1,J2MID_EFb_END1,J2MID_CDb_END1,J2MID_ABb_END1,W1END3,SS4END1,E1END3,NN4END1,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_W6BEG0 (
    .A0(W6BEG0_input[0]),
    .A1(W6BEG0_input[1]),
    .A2(W6BEG0_input[2]),
    .A3(W6BEG0_input[3]),
    .A4(W6BEG0_input[4]),
    .A5(W6BEG0_input[5]),
    .A6(W6BEG0_input[6]),
    .A7(W6BEG0_input[7]),
    .A8(W6BEG0_input[8]),
    .A9(W6BEG0_input[9]),
    .A10(W6BEG0_input[10]),
    .A11(W6BEG0_input[11]),
    .A12(W6BEG0_input[12]),
    .A13(W6BEG0_input[13]),
    .A14(W6BEG0_input[14]),
    .A15(W6BEG0_input[15]),
    .S0(ConfigBits[120+0]),
    .S0N(ConfigBits_N[120+0]),
    .S1(ConfigBits[120+1]),
    .S1N(ConfigBits_N[120+1]),
    .S2(ConfigBits[120+2]),
    .S2N(ConfigBits_N[120+2]),
    .S3(ConfigBits[120+3]),
    .S3N(ConfigBits_N[120+3]),
    .X(W6BEG0)
);

 //switch matrix multiplexer W6BEG1 MUX-16
assign W6BEG1_input = {J2MID_GHa_END2,J2MID_EFa_END2,J2MID_CDa_END2,J2MID_ABa_END2,W1END2,SS4END2,E1END2,NN4END2,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_W6BEG1 (
    .A0(W6BEG1_input[0]),
    .A1(W6BEG1_input[1]),
    .A2(W6BEG1_input[2]),
    .A3(W6BEG1_input[3]),
    .A4(W6BEG1_input[4]),
    .A5(W6BEG1_input[5]),
    .A6(W6BEG1_input[6]),
    .A7(W6BEG1_input[7]),
    .A8(W6BEG1_input[8]),
    .A9(W6BEG1_input[9]),
    .A10(W6BEG1_input[10]),
    .A11(W6BEG1_input[11]),
    .A12(W6BEG1_input[12]),
    .A13(W6BEG1_input[13]),
    .A14(W6BEG1_input[14]),
    .A15(W6BEG1_input[15]),
    .S0(ConfigBits[124+0]),
    .S0N(ConfigBits_N[124+0]),
    .S1(ConfigBits[124+1]),
    .S1N(ConfigBits_N[124+1]),
    .S2(ConfigBits[124+2]),
    .S2N(ConfigBits_N[124+2]),
    .S3(ConfigBits[124+3]),
    .S3N(ConfigBits_N[124+3]),
    .X(W6BEG1)
);

 //switch matrix multiplexer J2MID_ABa_BEG0 MUX-4
assign J2MID_ABa_BEG0_input = {JN2END3,W2MID6,S2MID6,N2MID6};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG0 (
    .A0(J2MID_ABa_BEG0_input[0]),
    .A1(J2MID_ABa_BEG0_input[1]),
    .A2(J2MID_ABa_BEG0_input[2]),
    .A3(J2MID_ABa_BEG0_input[3]),
    .S0(ConfigBits[128+0]),
    .S0N(ConfigBits_N[128+0]),
    .S1(ConfigBits[128+1]),
    .S1N(ConfigBits_N[128+1]),
    .X(J2MID_ABa_BEG0)
);

 //switch matrix multiplexer J2MID_ABa_BEG1 MUX-4
assign J2MID_ABa_BEG1_input = {JE2END3,W2MID2,S2MID2,E2MID2};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG1 (
    .A0(J2MID_ABa_BEG1_input[0]),
    .A1(J2MID_ABa_BEG1_input[1]),
    .A2(J2MID_ABa_BEG1_input[2]),
    .A3(J2MID_ABa_BEG1_input[3]),
    .S0(ConfigBits[130+0]),
    .S0N(ConfigBits_N[130+0]),
    .S1(ConfigBits[130+1]),
    .S1N(ConfigBits_N[130+1]),
    .X(J2MID_ABa_BEG1)
);

 //switch matrix multiplexer J2MID_ABa_BEG2 MUX-4
assign J2MID_ABa_BEG2_input = {JS2END3,W2MID4,E2MID4,N2MID4};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG2 (
    .A0(J2MID_ABa_BEG2_input[0]),
    .A1(J2MID_ABa_BEG2_input[1]),
    .A2(J2MID_ABa_BEG2_input[2]),
    .A3(J2MID_ABa_BEG2_input[3]),
    .S0(ConfigBits[132+0]),
    .S0N(ConfigBits_N[132+0]),
    .S1(ConfigBits[132+1]),
    .S1N(ConfigBits_N[132+1]),
    .X(J2MID_ABa_BEG2)
);

 //switch matrix multiplexer J2MID_ABa_BEG3 MUX-4
assign J2MID_ABa_BEG3_input = {JW2END3,S2MID0,E2MID0,N2MID0};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG3 (
    .A0(J2MID_ABa_BEG3_input[0]),
    .A1(J2MID_ABa_BEG3_input[1]),
    .A2(J2MID_ABa_BEG3_input[2]),
    .A3(J2MID_ABa_BEG3_input[3]),
    .S0(ConfigBits[134+0]),
    .S0N(ConfigBits_N[134+0]),
    .S1(ConfigBits[134+1]),
    .S1N(ConfigBits_N[134+1]),
    .X(J2MID_ABa_BEG3)
);

 //switch matrix multiplexer J2MID_CDa_BEG0 MUX-4
assign J2MID_CDa_BEG0_input = {JN2END4,W2MID6,S2MID6,E2MID6};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG0 (
    .A0(J2MID_CDa_BEG0_input[0]),
    .A1(J2MID_CDa_BEG0_input[1]),
    .A2(J2MID_CDa_BEG0_input[2]),
    .A3(J2MID_CDa_BEG0_input[3]),
    .S0(ConfigBits[136+0]),
    .S0N(ConfigBits_N[136+0]),
    .S1(ConfigBits[136+1]),
    .S1N(ConfigBits_N[136+1]),
    .X(J2MID_CDa_BEG0)
);

 //switch matrix multiplexer J2MID_CDa_BEG1 MUX-4
assign J2MID_CDa_BEG1_input = {JE2END4,W2MID2,E2MID2,N2MID2};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG1 (
    .A0(J2MID_CDa_BEG1_input[0]),
    .A1(J2MID_CDa_BEG1_input[1]),
    .A2(J2MID_CDa_BEG1_input[2]),
    .A3(J2MID_CDa_BEG1_input[3]),
    .S0(ConfigBits[138+0]),
    .S0N(ConfigBits_N[138+0]),
    .S1(ConfigBits[138+1]),
    .S1N(ConfigBits_N[138+1]),
    .X(J2MID_CDa_BEG1)
);

 //switch matrix multiplexer J2MID_CDa_BEG2 MUX-4
assign J2MID_CDa_BEG2_input = {JS2END4,S2MID4,E2MID4,N2MID4};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG2 (
    .A0(J2MID_CDa_BEG2_input[0]),
    .A1(J2MID_CDa_BEG2_input[1]),
    .A2(J2MID_CDa_BEG2_input[2]),
    .A3(J2MID_CDa_BEG2_input[3]),
    .S0(ConfigBits[140+0]),
    .S0N(ConfigBits_N[140+0]),
    .S1(ConfigBits[140+1]),
    .S1N(ConfigBits_N[140+1]),
    .X(J2MID_CDa_BEG2)
);

 //switch matrix multiplexer J2MID_CDa_BEG3 MUX-4
assign J2MID_CDa_BEG3_input = {JW2END4,W2MID0,S2MID0,N2MID0};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG3 (
    .A0(J2MID_CDa_BEG3_input[0]),
    .A1(J2MID_CDa_BEG3_input[1]),
    .A2(J2MID_CDa_BEG3_input[2]),
    .A3(J2MID_CDa_BEG3_input[3]),
    .S0(ConfigBits[142+0]),
    .S0N(ConfigBits_N[142+0]),
    .S1(ConfigBits[142+1]),
    .S1N(ConfigBits_N[142+1]),
    .X(J2MID_CDa_BEG3)
);

 //switch matrix multiplexer J2MID_EFa_BEG0 MUX-4
assign J2MID_EFa_BEG0_input = {JN2END5,W2MID6,E2MID6,N2MID6};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG0 (
    .A0(J2MID_EFa_BEG0_input[0]),
    .A1(J2MID_EFa_BEG0_input[1]),
    .A2(J2MID_EFa_BEG0_input[2]),
    .A3(J2MID_EFa_BEG0_input[3]),
    .S0(ConfigBits[144+0]),
    .S0N(ConfigBits_N[144+0]),
    .S1(ConfigBits[144+1]),
    .S1N(ConfigBits_N[144+1]),
    .X(J2MID_EFa_BEG0)
);

 //switch matrix multiplexer J2MID_EFa_BEG1 MUX-4
assign J2MID_EFa_BEG1_input = {JE2END5,S2MID2,E2MID2,N2MID2};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG1 (
    .A0(J2MID_EFa_BEG1_input[0]),
    .A1(J2MID_EFa_BEG1_input[1]),
    .A2(J2MID_EFa_BEG1_input[2]),
    .A3(J2MID_EFa_BEG1_input[3]),
    .S0(ConfigBits[146+0]),
    .S0N(ConfigBits_N[146+0]),
    .S1(ConfigBits[146+1]),
    .S1N(ConfigBits_N[146+1]),
    .X(J2MID_EFa_BEG1)
);

 //switch matrix multiplexer J2MID_EFa_BEG2 MUX-4
assign J2MID_EFa_BEG2_input = {JS2END5,W2MID4,S2MID4,N2MID4};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG2 (
    .A0(J2MID_EFa_BEG2_input[0]),
    .A1(J2MID_EFa_BEG2_input[1]),
    .A2(J2MID_EFa_BEG2_input[2]),
    .A3(J2MID_EFa_BEG2_input[3]),
    .S0(ConfigBits[148+0]),
    .S0N(ConfigBits_N[148+0]),
    .S1(ConfigBits[148+1]),
    .S1N(ConfigBits_N[148+1]),
    .X(J2MID_EFa_BEG2)
);

 //switch matrix multiplexer J2MID_EFa_BEG3 MUX-4
assign J2MID_EFa_BEG3_input = {JW2END5,W2MID0,S2MID0,E2MID0};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG3 (
    .A0(J2MID_EFa_BEG3_input[0]),
    .A1(J2MID_EFa_BEG3_input[1]),
    .A2(J2MID_EFa_BEG3_input[2]),
    .A3(J2MID_EFa_BEG3_input[3]),
    .S0(ConfigBits[150+0]),
    .S0N(ConfigBits_N[150+0]),
    .S1(ConfigBits[150+1]),
    .S1N(ConfigBits_N[150+1]),
    .X(J2MID_EFa_BEG3)
);

 //switch matrix multiplexer J2MID_GHa_BEG0 MUX-4
assign J2MID_GHa_BEG0_input = {JN2END6,S2MID6,E2MID6,N2MID6};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG0 (
    .A0(J2MID_GHa_BEG0_input[0]),
    .A1(J2MID_GHa_BEG0_input[1]),
    .A2(J2MID_GHa_BEG0_input[2]),
    .A3(J2MID_GHa_BEG0_input[3]),
    .S0(ConfigBits[152+0]),
    .S0N(ConfigBits_N[152+0]),
    .S1(ConfigBits[152+1]),
    .S1N(ConfigBits_N[152+1]),
    .X(J2MID_GHa_BEG0)
);

 //switch matrix multiplexer J2MID_GHa_BEG1 MUX-4
assign J2MID_GHa_BEG1_input = {JE2END6,W2MID2,S2MID2,N2MID2};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG1 (
    .A0(J2MID_GHa_BEG1_input[0]),
    .A1(J2MID_GHa_BEG1_input[1]),
    .A2(J2MID_GHa_BEG1_input[2]),
    .A3(J2MID_GHa_BEG1_input[3]),
    .S0(ConfigBits[154+0]),
    .S0N(ConfigBits_N[154+0]),
    .S1(ConfigBits[154+1]),
    .S1N(ConfigBits_N[154+1]),
    .X(J2MID_GHa_BEG1)
);

 //switch matrix multiplexer J2MID_GHa_BEG2 MUX-4
assign J2MID_GHa_BEG2_input = {JS2END6,W2MID4,S2MID4,E2MID4};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG2 (
    .A0(J2MID_GHa_BEG2_input[0]),
    .A1(J2MID_GHa_BEG2_input[1]),
    .A2(J2MID_GHa_BEG2_input[2]),
    .A3(J2MID_GHa_BEG2_input[3]),
    .S0(ConfigBits[156+0]),
    .S0N(ConfigBits_N[156+0]),
    .S1(ConfigBits[156+1]),
    .S1N(ConfigBits_N[156+1]),
    .X(J2MID_GHa_BEG2)
);

 //switch matrix multiplexer J2MID_GHa_BEG3 MUX-4
assign J2MID_GHa_BEG3_input = {JW2END6,W2MID0,E2MID0,N2MID0};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG3 (
    .A0(J2MID_GHa_BEG3_input[0]),
    .A1(J2MID_GHa_BEG3_input[1]),
    .A2(J2MID_GHa_BEG3_input[2]),
    .A3(J2MID_GHa_BEG3_input[3]),
    .S0(ConfigBits[158+0]),
    .S0N(ConfigBits_N[158+0]),
    .S1(ConfigBits[158+1]),
    .S1N(ConfigBits_N[158+1]),
    .X(J2MID_GHa_BEG3)
);

 //switch matrix multiplexer J2MID_ABb_BEG0 MUX-4
assign J2MID_ABb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG0 (
    .A0(J2MID_ABb_BEG0_input[0]),
    .A1(J2MID_ABb_BEG0_input[1]),
    .A2(J2MID_ABb_BEG0_input[2]),
    .A3(J2MID_ABb_BEG0_input[3]),
    .S0(ConfigBits[160+0]),
    .S0N(ConfigBits_N[160+0]),
    .S1(ConfigBits[160+1]),
    .S1N(ConfigBits_N[160+1]),
    .X(J2MID_ABb_BEG0)
);

 //switch matrix multiplexer J2MID_ABb_BEG1 MUX-4
assign J2MID_ABb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG1 (
    .A0(J2MID_ABb_BEG1_input[0]),
    .A1(J2MID_ABb_BEG1_input[1]),
    .A2(J2MID_ABb_BEG1_input[2]),
    .A3(J2MID_ABb_BEG1_input[3]),
    .S0(ConfigBits[162+0]),
    .S0N(ConfigBits_N[162+0]),
    .S1(ConfigBits[162+1]),
    .S1N(ConfigBits_N[162+1]),
    .X(J2MID_ABb_BEG1)
);

 //switch matrix multiplexer J2MID_ABb_BEG2 MUX-4
assign J2MID_ABb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG2 (
    .A0(J2MID_ABb_BEG2_input[0]),
    .A1(J2MID_ABb_BEG2_input[1]),
    .A2(J2MID_ABb_BEG2_input[2]),
    .A3(J2MID_ABb_BEG2_input[3]),
    .S0(ConfigBits[164+0]),
    .S0N(ConfigBits_N[164+0]),
    .S1(ConfigBits[164+1]),
    .S1N(ConfigBits_N[164+1]),
    .X(J2MID_ABb_BEG2)
);

 //switch matrix multiplexer J2MID_ABb_BEG3 MUX-4
assign J2MID_ABb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG3 (
    .A0(J2MID_ABb_BEG3_input[0]),
    .A1(J2MID_ABb_BEG3_input[1]),
    .A2(J2MID_ABb_BEG3_input[2]),
    .A3(J2MID_ABb_BEG3_input[3]),
    .S0(ConfigBits[166+0]),
    .S0N(ConfigBits_N[166+0]),
    .S1(ConfigBits[166+1]),
    .S1N(ConfigBits_N[166+1]),
    .X(J2MID_ABb_BEG3)
);

 //switch matrix multiplexer J2MID_CDb_BEG0 MUX-4
assign J2MID_CDb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG0 (
    .A0(J2MID_CDb_BEG0_input[0]),
    .A1(J2MID_CDb_BEG0_input[1]),
    .A2(J2MID_CDb_BEG0_input[2]),
    .A3(J2MID_CDb_BEG0_input[3]),
    .S0(ConfigBits[168+0]),
    .S0N(ConfigBits_N[168+0]),
    .S1(ConfigBits[168+1]),
    .S1N(ConfigBits_N[168+1]),
    .X(J2MID_CDb_BEG0)
);

 //switch matrix multiplexer J2MID_CDb_BEG1 MUX-4
assign J2MID_CDb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG1 (
    .A0(J2MID_CDb_BEG1_input[0]),
    .A1(J2MID_CDb_BEG1_input[1]),
    .A2(J2MID_CDb_BEG1_input[2]),
    .A3(J2MID_CDb_BEG1_input[3]),
    .S0(ConfigBits[170+0]),
    .S0N(ConfigBits_N[170+0]),
    .S1(ConfigBits[170+1]),
    .S1N(ConfigBits_N[170+1]),
    .X(J2MID_CDb_BEG1)
);

 //switch matrix multiplexer J2MID_CDb_BEG2 MUX-4
assign J2MID_CDb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG2 (
    .A0(J2MID_CDb_BEG2_input[0]),
    .A1(J2MID_CDb_BEG2_input[1]),
    .A2(J2MID_CDb_BEG2_input[2]),
    .A3(J2MID_CDb_BEG2_input[3]),
    .S0(ConfigBits[172+0]),
    .S0N(ConfigBits_N[172+0]),
    .S1(ConfigBits[172+1]),
    .S1N(ConfigBits_N[172+1]),
    .X(J2MID_CDb_BEG2)
);

 //switch matrix multiplexer J2MID_CDb_BEG3 MUX-4
assign J2MID_CDb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG3 (
    .A0(J2MID_CDb_BEG3_input[0]),
    .A1(J2MID_CDb_BEG3_input[1]),
    .A2(J2MID_CDb_BEG3_input[2]),
    .A3(J2MID_CDb_BEG3_input[3]),
    .S0(ConfigBits[174+0]),
    .S0N(ConfigBits_N[174+0]),
    .S1(ConfigBits[174+1]),
    .S1N(ConfigBits_N[174+1]),
    .X(J2MID_CDb_BEG3)
);

 //switch matrix multiplexer J2MID_EFb_BEG0 MUX-4
assign J2MID_EFb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG0 (
    .A0(J2MID_EFb_BEG0_input[0]),
    .A1(J2MID_EFb_BEG0_input[1]),
    .A2(J2MID_EFb_BEG0_input[2]),
    .A3(J2MID_EFb_BEG0_input[3]),
    .S0(ConfigBits[176+0]),
    .S0N(ConfigBits_N[176+0]),
    .S1(ConfigBits[176+1]),
    .S1N(ConfigBits_N[176+1]),
    .X(J2MID_EFb_BEG0)
);

 //switch matrix multiplexer J2MID_EFb_BEG1 MUX-4
assign J2MID_EFb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG1 (
    .A0(J2MID_EFb_BEG1_input[0]),
    .A1(J2MID_EFb_BEG1_input[1]),
    .A2(J2MID_EFb_BEG1_input[2]),
    .A3(J2MID_EFb_BEG1_input[3]),
    .S0(ConfigBits[178+0]),
    .S0N(ConfigBits_N[178+0]),
    .S1(ConfigBits[178+1]),
    .S1N(ConfigBits_N[178+1]),
    .X(J2MID_EFb_BEG1)
);

 //switch matrix multiplexer J2MID_EFb_BEG2 MUX-4
assign J2MID_EFb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG2 (
    .A0(J2MID_EFb_BEG2_input[0]),
    .A1(J2MID_EFb_BEG2_input[1]),
    .A2(J2MID_EFb_BEG2_input[2]),
    .A3(J2MID_EFb_BEG2_input[3]),
    .S0(ConfigBits[180+0]),
    .S0N(ConfigBits_N[180+0]),
    .S1(ConfigBits[180+1]),
    .S1N(ConfigBits_N[180+1]),
    .X(J2MID_EFb_BEG2)
);

 //switch matrix multiplexer J2MID_EFb_BEG3 MUX-4
assign J2MID_EFb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG3 (
    .A0(J2MID_EFb_BEG3_input[0]),
    .A1(J2MID_EFb_BEG3_input[1]),
    .A2(J2MID_EFb_BEG3_input[2]),
    .A3(J2MID_EFb_BEG3_input[3]),
    .S0(ConfigBits[182+0]),
    .S0N(ConfigBits_N[182+0]),
    .S1(ConfigBits[182+1]),
    .S1N(ConfigBits_N[182+1]),
    .X(J2MID_EFb_BEG3)
);

 //switch matrix multiplexer J2MID_GHb_BEG0 MUX-4
assign J2MID_GHb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG0 (
    .A0(J2MID_GHb_BEG0_input[0]),
    .A1(J2MID_GHb_BEG0_input[1]),
    .A2(J2MID_GHb_BEG0_input[2]),
    .A3(J2MID_GHb_BEG0_input[3]),
    .S0(ConfigBits[184+0]),
    .S0N(ConfigBits_N[184+0]),
    .S1(ConfigBits[184+1]),
    .S1N(ConfigBits_N[184+1]),
    .X(J2MID_GHb_BEG0)
);

 //switch matrix multiplexer J2MID_GHb_BEG1 MUX-4
assign J2MID_GHb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG1 (
    .A0(J2MID_GHb_BEG1_input[0]),
    .A1(J2MID_GHb_BEG1_input[1]),
    .A2(J2MID_GHb_BEG1_input[2]),
    .A3(J2MID_GHb_BEG1_input[3]),
    .S0(ConfigBits[186+0]),
    .S0N(ConfigBits_N[186+0]),
    .S1(ConfigBits[186+1]),
    .S1N(ConfigBits_N[186+1]),
    .X(J2MID_GHb_BEG1)
);

 //switch matrix multiplexer J2MID_GHb_BEG2 MUX-4
assign J2MID_GHb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG2 (
    .A0(J2MID_GHb_BEG2_input[0]),
    .A1(J2MID_GHb_BEG2_input[1]),
    .A2(J2MID_GHb_BEG2_input[2]),
    .A3(J2MID_GHb_BEG2_input[3]),
    .S0(ConfigBits[188+0]),
    .S0N(ConfigBits_N[188+0]),
    .S1(ConfigBits[188+1]),
    .S1N(ConfigBits_N[188+1]),
    .X(J2MID_GHb_BEG2)
);

 //switch matrix multiplexer J2MID_GHb_BEG3 MUX-4
assign J2MID_GHb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG3 (
    .A0(J2MID_GHb_BEG3_input[0]),
    .A1(J2MID_GHb_BEG3_input[1]),
    .A2(J2MID_GHb_BEG3_input[2]),
    .A3(J2MID_GHb_BEG3_input[3]),
    .S0(ConfigBits[190+0]),
    .S0N(ConfigBits_N[190+0]),
    .S1(ConfigBits[190+1]),
    .S1N(ConfigBits_N[190+1]),
    .X(J2MID_GHb_BEG3)
);

 //switch matrix multiplexer J2END_AB_BEG0 MUX-4
assign J2END_AB_BEG0_input = {W2END6,SS4END3,E2END6,N2END6};
cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG0 (
    .A0(J2END_AB_BEG0_input[0]),
    .A1(J2END_AB_BEG0_input[1]),
    .A2(J2END_AB_BEG0_input[2]),
    .A3(J2END_AB_BEG0_input[3]),
    .S0(ConfigBits[192+0]),
    .S0N(ConfigBits_N[192+0]),
    .S1(ConfigBits[192+1]),
    .S1N(ConfigBits_N[192+1]),
    .X(J2END_AB_BEG0)
);

 //switch matrix multiplexer J2END_AB_BEG1 MUX-4
assign J2END_AB_BEG1_input = {W2END2,S2END2,E2END2,NN4END0};
cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG1 (
    .A0(J2END_AB_BEG1_input[0]),
    .A1(J2END_AB_BEG1_input[1]),
    .A2(J2END_AB_BEG1_input[2]),
    .A3(J2END_AB_BEG1_input[3]),
    .S0(ConfigBits[194+0]),
    .S0N(ConfigBits_N[194+0]),
    .S1(ConfigBits[194+1]),
    .S1N(ConfigBits_N[194+1]),
    .X(J2END_AB_BEG1)
);

 //switch matrix multiplexer J2END_AB_BEG2 MUX-4
assign J2END_AB_BEG2_input = {W2END4,S2END4,EE4END0,N2END4};
cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG2 (
    .A0(J2END_AB_BEG2_input[0]),
    .A1(J2END_AB_BEG2_input[1]),
    .A2(J2END_AB_BEG2_input[2]),
    .A3(J2END_AB_BEG2_input[3]),
    .S0(ConfigBits[196+0]),
    .S0N(ConfigBits_N[196+0]),
    .S1(ConfigBits[196+1]),
    .S1N(ConfigBits_N[196+1]),
    .X(J2END_AB_BEG2)
);

 //switch matrix multiplexer J2END_AB_BEG3 MUX-4
assign J2END_AB_BEG3_input = {WW4END3,S2END0,E2END0,N2END0};
cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG3 (
    .A0(J2END_AB_BEG3_input[0]),
    .A1(J2END_AB_BEG3_input[1]),
    .A2(J2END_AB_BEG3_input[2]),
    .A3(J2END_AB_BEG3_input[3]),
    .S0(ConfigBits[198+0]),
    .S0N(ConfigBits_N[198+0]),
    .S1(ConfigBits[198+1]),
    .S1N(ConfigBits_N[198+1]),
    .X(J2END_AB_BEG3)
);

 //switch matrix multiplexer J2END_CD_BEG0 MUX-4
assign J2END_CD_BEG0_input = {W2END6,S2END6,E2END6,NN4END3};
cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG0 (
    .A0(J2END_CD_BEG0_input[0]),
    .A1(J2END_CD_BEG0_input[1]),
    .A2(J2END_CD_BEG0_input[2]),
    .A3(J2END_CD_BEG0_input[3]),
    .S0(ConfigBits[200+0]),
    .S0N(ConfigBits_N[200+0]),
    .S1(ConfigBits[200+1]),
    .S1N(ConfigBits_N[200+1]),
    .X(J2END_CD_BEG0)
);

 //switch matrix multiplexer J2END_CD_BEG1 MUX-4
assign J2END_CD_BEG1_input = {WW4END2,S2END2,E2END2,N2END2};
cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG1 (
    .A0(J2END_CD_BEG1_input[0]),
    .A1(J2END_CD_BEG1_input[1]),
    .A2(J2END_CD_BEG1_input[2]),
    .A3(J2END_CD_BEG1_input[3]),
    .S0(ConfigBits[202+0]),
    .S0N(ConfigBits_N[202+0]),
    .S1(ConfigBits[202+1]),
    .S1N(ConfigBits_N[202+1]),
    .X(J2END_CD_BEG1)
);

 //switch matrix multiplexer J2END_CD_BEG2 MUX-4
assign J2END_CD_BEG2_input = {W2END4,SS4END2,E2END4,N2END4};
cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG2 (
    .A0(J2END_CD_BEG2_input[0]),
    .A1(J2END_CD_BEG2_input[1]),
    .A2(J2END_CD_BEG2_input[2]),
    .A3(J2END_CD_BEG2_input[3]),
    .S0(ConfigBits[204+0]),
    .S0N(ConfigBits_N[204+0]),
    .S1(ConfigBits[204+1]),
    .S1N(ConfigBits_N[204+1]),
    .X(J2END_CD_BEG2)
);

 //switch matrix multiplexer J2END_CD_BEG3 MUX-4
assign J2END_CD_BEG3_input = {W2END0,S2END0,EE4END1,N2END0};
cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG3 (
    .A0(J2END_CD_BEG3_input[0]),
    .A1(J2END_CD_BEG3_input[1]),
    .A2(J2END_CD_BEG3_input[2]),
    .A3(J2END_CD_BEG3_input[3]),
    .S0(ConfigBits[206+0]),
    .S0N(ConfigBits_N[206+0]),
    .S1(ConfigBits[206+1]),
    .S1N(ConfigBits_N[206+1]),
    .X(J2END_CD_BEG3)
);

 //switch matrix multiplexer J2END_EF_BEG0 MUX-4
assign J2END_EF_BEG0_input = {W2END7,S2END7,EE4END2,N2END7};
cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG0 (
    .A0(J2END_EF_BEG0_input[0]),
    .A1(J2END_EF_BEG0_input[1]),
    .A2(J2END_EF_BEG0_input[2]),
    .A3(J2END_EF_BEG0_input[3]),
    .S0(ConfigBits[208+0]),
    .S0N(ConfigBits_N[208+0]),
    .S1(ConfigBits[208+1]),
    .S1N(ConfigBits_N[208+1]),
    .X(J2END_EF_BEG0)
);

 //switch matrix multiplexer J2END_EF_BEG1 MUX-4
assign J2END_EF_BEG1_input = {WW4END1,S2END3,E2END3,N2END3};
cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG1 (
    .A0(J2END_EF_BEG1_input[0]),
    .A1(J2END_EF_BEG1_input[1]),
    .A2(J2END_EF_BEG1_input[2]),
    .A3(J2END_EF_BEG1_input[3]),
    .S0(ConfigBits[210+0]),
    .S0N(ConfigBits_N[210+0]),
    .S1(ConfigBits[210+1]),
    .S1N(ConfigBits_N[210+1]),
    .X(J2END_EF_BEG1)
);

 //switch matrix multiplexer J2END_EF_BEG2 MUX-4
assign J2END_EF_BEG2_input = {W2END5,SS4END1,E2END5,N2END5};
cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG2 (
    .A0(J2END_EF_BEG2_input[0]),
    .A1(J2END_EF_BEG2_input[1]),
    .A2(J2END_EF_BEG2_input[2]),
    .A3(J2END_EF_BEG2_input[3]),
    .S0(ConfigBits[212+0]),
    .S0N(ConfigBits_N[212+0]),
    .S1(ConfigBits[212+1]),
    .S1N(ConfigBits_N[212+1]),
    .X(J2END_EF_BEG2)
);

 //switch matrix multiplexer J2END_EF_BEG3 MUX-4
assign J2END_EF_BEG3_input = {W2END1,S2END1,E2END1,NN4END2};
cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG3 (
    .A0(J2END_EF_BEG3_input[0]),
    .A1(J2END_EF_BEG3_input[1]),
    .A2(J2END_EF_BEG3_input[2]),
    .A3(J2END_EF_BEG3_input[3]),
    .S0(ConfigBits[214+0]),
    .S0N(ConfigBits_N[214+0]),
    .S1(ConfigBits[214+1]),
    .S1N(ConfigBits_N[214+1]),
    .X(J2END_EF_BEG3)
);

 //switch matrix multiplexer J2END_GH_BEG0 MUX-4
assign J2END_GH_BEG0_input = {WW4END0,S2END7,E2END7,N2END7};
cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG0 (
    .A0(J2END_GH_BEG0_input[0]),
    .A1(J2END_GH_BEG0_input[1]),
    .A2(J2END_GH_BEG0_input[2]),
    .A3(J2END_GH_BEG0_input[3]),
    .S0(ConfigBits[216+0]),
    .S0N(ConfigBits_N[216+0]),
    .S1(ConfigBits[216+1]),
    .S1N(ConfigBits_N[216+1]),
    .X(J2END_GH_BEG0)
);

 //switch matrix multiplexer J2END_GH_BEG1 MUX-4
assign J2END_GH_BEG1_input = {W2END3,SS4END0,E2END3,N2END3};
cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG1 (
    .A0(J2END_GH_BEG1_input[0]),
    .A1(J2END_GH_BEG1_input[1]),
    .A2(J2END_GH_BEG1_input[2]),
    .A3(J2END_GH_BEG1_input[3]),
    .S0(ConfigBits[218+0]),
    .S0N(ConfigBits_N[218+0]),
    .S1(ConfigBits[218+1]),
    .S1N(ConfigBits_N[218+1]),
    .X(J2END_GH_BEG1)
);

 //switch matrix multiplexer J2END_GH_BEG2 MUX-4
assign J2END_GH_BEG2_input = {W2END5,S2END5,E2END5,NN4END1};
cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG2 (
    .A0(J2END_GH_BEG2_input[0]),
    .A1(J2END_GH_BEG2_input[1]),
    .A2(J2END_GH_BEG2_input[2]),
    .A3(J2END_GH_BEG2_input[3]),
    .S0(ConfigBits[220+0]),
    .S0N(ConfigBits_N[220+0]),
    .S1(ConfigBits[220+1]),
    .S1N(ConfigBits_N[220+1]),
    .X(J2END_GH_BEG2)
);

 //switch matrix multiplexer J2END_GH_BEG3 MUX-4
assign J2END_GH_BEG3_input = {W2END1,S2END1,EE4END3,N2END1};
cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG3 (
    .A0(J2END_GH_BEG3_input[0]),
    .A1(J2END_GH_BEG3_input[1]),
    .A2(J2END_GH_BEG3_input[2]),
    .A3(J2END_GH_BEG3_input[3]),
    .S0(ConfigBits[222+0]),
    .S0N(ConfigBits_N[222+0]),
    .S1(ConfigBits[222+1]),
    .S1N(ConfigBits_N[222+1]),
    .X(J2END_GH_BEG3)
);

 //switch matrix multiplexer JN2BEG0 MUX-16
assign JN2BEG0_input = {W6END1,W2END1,S2END1,E6END1,EE4END0,E2END1,E1END3,N4END1,N2END1,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG0 (
    .A0(JN2BEG0_input[0]),
    .A1(JN2BEG0_input[1]),
    .A2(JN2BEG0_input[2]),
    .A3(JN2BEG0_input[3]),
    .A4(JN2BEG0_input[4]),
    .A5(JN2BEG0_input[5]),
    .A6(JN2BEG0_input[6]),
    .A7(JN2BEG0_input[7]),
    .A8(JN2BEG0_input[8]),
    .A9(JN2BEG0_input[9]),
    .A10(JN2BEG0_input[10]),
    .A11(JN2BEG0_input[11]),
    .A12(JN2BEG0_input[12]),
    .A13(JN2BEG0_input[13]),
    .A14(JN2BEG0_input[14]),
    .A15(JN2BEG0_input[15]),
    .S0(ConfigBits[224+0]),
    .S0N(ConfigBits_N[224+0]),
    .S1(ConfigBits[224+1]),
    .S1N(ConfigBits_N[224+1]),
    .S2(ConfigBits[224+2]),
    .S2N(ConfigBits_N[224+2]),
    .S3(ConfigBits[224+3]),
    .S3N(ConfigBits_N[224+3]),
    .X(JN2BEG0)
);

 //switch matrix multiplexer JN2BEG1 MUX-16
assign JN2BEG1_input = {W6END0,W2END2,S2END2,E6END0,EE4END1,E2END2,E1END0,N4END2,N2END2,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG1 (
    .A0(JN2BEG1_input[0]),
    .A1(JN2BEG1_input[1]),
    .A2(JN2BEG1_input[2]),
    .A3(JN2BEG1_input[3]),
    .A4(JN2BEG1_input[4]),
    .A5(JN2BEG1_input[5]),
    .A6(JN2BEG1_input[6]),
    .A7(JN2BEG1_input[7]),
    .A8(JN2BEG1_input[8]),
    .A9(JN2BEG1_input[9]),
    .A10(JN2BEG1_input[10]),
    .A11(JN2BEG1_input[11]),
    .A12(JN2BEG1_input[12]),
    .A13(JN2BEG1_input[13]),
    .A14(JN2BEG1_input[14]),
    .A15(JN2BEG1_input[15]),
    .S0(ConfigBits[228+0]),
    .S0N(ConfigBits_N[228+0]),
    .S1(ConfigBits[228+1]),
    .S1N(ConfigBits_N[228+1]),
    .S2(ConfigBits[228+2]),
    .S2N(ConfigBits_N[228+2]),
    .S3(ConfigBits[228+3]),
    .S3N(ConfigBits_N[228+3]),
    .X(JN2BEG1)
);

 //switch matrix multiplexer JN2BEG2 MUX-16
assign JN2BEG2_input = {W6END1,WW4END2,W2END3,S2END3,E6END1,E2END3,E1END1,N4END3,N2END3,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG2 (
    .A0(JN2BEG2_input[0]),
    .A1(JN2BEG2_input[1]),
    .A2(JN2BEG2_input[2]),
    .A3(JN2BEG2_input[3]),
    .A4(JN2BEG2_input[4]),
    .A5(JN2BEG2_input[5]),
    .A6(JN2BEG2_input[6]),
    .A7(JN2BEG2_input[7]),
    .A8(JN2BEG2_input[8]),
    .A9(JN2BEG2_input[9]),
    .A10(JN2BEG2_input[10]),
    .A11(JN2BEG2_input[11]),
    .A12(JN2BEG2_input[12]),
    .A13(JN2BEG2_input[13]),
    .A14(JN2BEG2_input[14]),
    .A15(JN2BEG2_input[15]),
    .S0(ConfigBits[232+0]),
    .S0N(ConfigBits_N[232+0]),
    .S1(ConfigBits[232+1]),
    .S1N(ConfigBits_N[232+1]),
    .S2(ConfigBits[232+2]),
    .S2N(ConfigBits_N[232+2]),
    .S3(ConfigBits[232+3]),
    .S3N(ConfigBits_N[232+3]),
    .X(JN2BEG2)
);

 //switch matrix multiplexer JN2BEG3 MUX-16
assign JN2BEG3_input = {W6END0,WW4END3,W2END4,S2END4,E6END0,E2END4,E1END2,N4END0,N2END4,o_6to27,o_6to26,o_6to25,o_6to24,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG3 (
    .A0(JN2BEG3_input[0]),
    .A1(JN2BEG3_input[1]),
    .A2(JN2BEG3_input[2]),
    .A3(JN2BEG3_input[3]),
    .A4(JN2BEG3_input[4]),
    .A5(JN2BEG3_input[5]),
    .A6(JN2BEG3_input[6]),
    .A7(JN2BEG3_input[7]),
    .A8(JN2BEG3_input[8]),
    .A9(JN2BEG3_input[9]),
    .A10(JN2BEG3_input[10]),
    .A11(JN2BEG3_input[11]),
    .A12(JN2BEG3_input[12]),
    .A13(JN2BEG3_input[13]),
    .A14(JN2BEG3_input[14]),
    .A15(JN2BEG3_input[15]),
    .S0(ConfigBits[236+0]),
    .S0N(ConfigBits_N[236+0]),
    .S1(ConfigBits[236+1]),
    .S1N(ConfigBits_N[236+1]),
    .S2(ConfigBits[236+2]),
    .S2N(ConfigBits_N[236+2]),
    .S3(ConfigBits[236+3]),
    .S3N(ConfigBits_N[236+3]),
    .X(JN2BEG3)
);

 //switch matrix multiplexer JN2BEG4 MUX-16
assign JN2BEG4_input = {W1END3,W1END1,S2END5,S1END1,E2END5,E1END1,NN4END3,N2END5,N1END1,o_6to27,o_6to26,o_6to25,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG4 (
    .A0(JN2BEG4_input[0]),
    .A1(JN2BEG4_input[1]),
    .A2(JN2BEG4_input[2]),
    .A3(JN2BEG4_input[3]),
    .A4(JN2BEG4_input[4]),
    .A5(JN2BEG4_input[5]),
    .A6(JN2BEG4_input[6]),
    .A7(JN2BEG4_input[7]),
    .A8(JN2BEG4_input[8]),
    .A9(JN2BEG4_input[9]),
    .A10(JN2BEG4_input[10]),
    .A11(JN2BEG4_input[11]),
    .A12(JN2BEG4_input[12]),
    .A13(JN2BEG4_input[13]),
    .A14(JN2BEG4_input[14]),
    .A15(JN2BEG4_input[15]),
    .S0(ConfigBits[240+0]),
    .S0N(ConfigBits_N[240+0]),
    .S1(ConfigBits[240+1]),
    .S1N(ConfigBits_N[240+1]),
    .S2(ConfigBits[240+2]),
    .S2N(ConfigBits_N[240+2]),
    .S3(ConfigBits[240+3]),
    .S3N(ConfigBits_N[240+3]),
    .X(JN2BEG4)
);

 //switch matrix multiplexer JN2BEG5 MUX-16
assign JN2BEG5_input = {W1END2,W1END0,S2END6,S1END2,E2END6,E1END2,NN4END2,N2END6,N1END2,o_6to27,o_6to26,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG5 (
    .A0(JN2BEG5_input[0]),
    .A1(JN2BEG5_input[1]),
    .A2(JN2BEG5_input[2]),
    .A3(JN2BEG5_input[3]),
    .A4(JN2BEG5_input[4]),
    .A5(JN2BEG5_input[5]),
    .A6(JN2BEG5_input[6]),
    .A7(JN2BEG5_input[7]),
    .A8(JN2BEG5_input[8]),
    .A9(JN2BEG5_input[9]),
    .A10(JN2BEG5_input[10]),
    .A11(JN2BEG5_input[11]),
    .A12(JN2BEG5_input[12]),
    .A13(JN2BEG5_input[13]),
    .A14(JN2BEG5_input[14]),
    .A15(JN2BEG5_input[15]),
    .S0(ConfigBits[244+0]),
    .S0N(ConfigBits_N[244+0]),
    .S1(ConfigBits[244+1]),
    .S1N(ConfigBits_N[244+1]),
    .S2(ConfigBits[244+2]),
    .S2N(ConfigBits_N[244+2]),
    .S3(ConfigBits[244+3]),
    .S3N(ConfigBits_N[244+3]),
    .X(JN2BEG5)
);

 //switch matrix multiplexer JN2BEG6 MUX-16
assign JN2BEG6_input = {W1END3,W1END1,S2END7,S1END3,E2END7,E1END3,NN4END1,N2END7,N1END3,o_6to27,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG6 (
    .A0(JN2BEG6_input[0]),
    .A1(JN2BEG6_input[1]),
    .A2(JN2BEG6_input[2]),
    .A3(JN2BEG6_input[3]),
    .A4(JN2BEG6_input[4]),
    .A5(JN2BEG6_input[5]),
    .A6(JN2BEG6_input[6]),
    .A7(JN2BEG6_input[7]),
    .A8(JN2BEG6_input[8]),
    .A9(JN2BEG6_input[9]),
    .A10(JN2BEG6_input[10]),
    .A11(JN2BEG6_input[11]),
    .A12(JN2BEG6_input[12]),
    .A13(JN2BEG6_input[13]),
    .A14(JN2BEG6_input[14]),
    .A15(JN2BEG6_input[15]),
    .S0(ConfigBits[248+0]),
    .S0N(ConfigBits_N[248+0]),
    .S1(ConfigBits[248+1]),
    .S1N(ConfigBits_N[248+1]),
    .S2(ConfigBits[248+2]),
    .S2N(ConfigBits_N[248+2]),
    .S3(ConfigBits[248+3]),
    .S3N(ConfigBits_N[248+3]),
    .X(JN2BEG6)
);

 //switch matrix multiplexer JN2BEG7 MUX-16
assign JN2BEG7_input = {W1END2,W1END0,S2END0,S1END0,E2END0,E1END0,NN4END0,N2END0,N1END0,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JN2BEG7 (
    .A0(JN2BEG7_input[0]),
    .A1(JN2BEG7_input[1]),
    .A2(JN2BEG7_input[2]),
    .A3(JN2BEG7_input[3]),
    .A4(JN2BEG7_input[4]),
    .A5(JN2BEG7_input[5]),
    .A6(JN2BEG7_input[6]),
    .A7(JN2BEG7_input[7]),
    .A8(JN2BEG7_input[8]),
    .A9(JN2BEG7_input[9]),
    .A10(JN2BEG7_input[10]),
    .A11(JN2BEG7_input[11]),
    .A12(JN2BEG7_input[12]),
    .A13(JN2BEG7_input[13]),
    .A14(JN2BEG7_input[14]),
    .A15(JN2BEG7_input[15]),
    .S0(ConfigBits[252+0]),
    .S0N(ConfigBits_N[252+0]),
    .S1(ConfigBits[252+1]),
    .S1N(ConfigBits_N[252+1]),
    .S2(ConfigBits[252+2]),
    .S2N(ConfigBits_N[252+2]),
    .S3(ConfigBits[252+3]),
    .S3N(ConfigBits_N[252+3]),
    .X(JN2BEG7)
);

 //switch matrix multiplexer JE2BEG0 MUX-16
assign JE2BEG0_input = {W6END1,W2END1,S2END1,E6END1,E2END1,NN4END0,N4END1,N2END1,N1END3,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG0 (
    .A0(JE2BEG0_input[0]),
    .A1(JE2BEG0_input[1]),
    .A2(JE2BEG0_input[2]),
    .A3(JE2BEG0_input[3]),
    .A4(JE2BEG0_input[4]),
    .A5(JE2BEG0_input[5]),
    .A6(JE2BEG0_input[6]),
    .A7(JE2BEG0_input[7]),
    .A8(JE2BEG0_input[8]),
    .A9(JE2BEG0_input[9]),
    .A10(JE2BEG0_input[10]),
    .A11(JE2BEG0_input[11]),
    .A12(JE2BEG0_input[12]),
    .A13(JE2BEG0_input[13]),
    .A14(JE2BEG0_input[14]),
    .A15(JE2BEG0_input[15]),
    .S0(ConfigBits[256+0]),
    .S0N(ConfigBits_N[256+0]),
    .S1(ConfigBits[256+1]),
    .S1N(ConfigBits_N[256+1]),
    .S2(ConfigBits[256+2]),
    .S2N(ConfigBits_N[256+2]),
    .S3(ConfigBits[256+3]),
    .S3N(ConfigBits_N[256+3]),
    .X(JE2BEG0)
);

 //switch matrix multiplexer JE2BEG1 MUX-16
assign JE2BEG1_input = {W6END0,W2END2,S2END2,E6END0,E2END2,NN4END1,N4END2,N2END2,N1END0,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG1 (
    .A0(JE2BEG1_input[0]),
    .A1(JE2BEG1_input[1]),
    .A2(JE2BEG1_input[2]),
    .A3(JE2BEG1_input[3]),
    .A4(JE2BEG1_input[4]),
    .A5(JE2BEG1_input[5]),
    .A6(JE2BEG1_input[6]),
    .A7(JE2BEG1_input[7]),
    .A8(JE2BEG1_input[8]),
    .A9(JE2BEG1_input[9]),
    .A10(JE2BEG1_input[10]),
    .A11(JE2BEG1_input[11]),
    .A12(JE2BEG1_input[12]),
    .A13(JE2BEG1_input[13]),
    .A14(JE2BEG1_input[14]),
    .A15(JE2BEG1_input[15]),
    .S0(ConfigBits[260+0]),
    .S0N(ConfigBits_N[260+0]),
    .S1(ConfigBits[260+1]),
    .S1N(ConfigBits_N[260+1]),
    .S2(ConfigBits[260+2]),
    .S2N(ConfigBits_N[260+2]),
    .S3(ConfigBits[260+3]),
    .S3N(ConfigBits_N[260+3]),
    .X(JE2BEG1)
);

 //switch matrix multiplexer JE2BEG2 MUX-16
assign JE2BEG2_input = {W6END1,W2END3,SS4END2,S2END3,E6END1,E2END3,N4END3,N2END3,N1END1,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG2 (
    .A0(JE2BEG2_input[0]),
    .A1(JE2BEG2_input[1]),
    .A2(JE2BEG2_input[2]),
    .A3(JE2BEG2_input[3]),
    .A4(JE2BEG2_input[4]),
    .A5(JE2BEG2_input[5]),
    .A6(JE2BEG2_input[6]),
    .A7(JE2BEG2_input[7]),
    .A8(JE2BEG2_input[8]),
    .A9(JE2BEG2_input[9]),
    .A10(JE2BEG2_input[10]),
    .A11(JE2BEG2_input[11]),
    .A12(JE2BEG2_input[12]),
    .A13(JE2BEG2_input[13]),
    .A14(JE2BEG2_input[14]),
    .A15(JE2BEG2_input[15]),
    .S0(ConfigBits[264+0]),
    .S0N(ConfigBits_N[264+0]),
    .S1(ConfigBits[264+1]),
    .S1N(ConfigBits_N[264+1]),
    .S2(ConfigBits[264+2]),
    .S2N(ConfigBits_N[264+2]),
    .S3(ConfigBits[264+3]),
    .S3N(ConfigBits_N[264+3]),
    .X(JE2BEG2)
);

 //switch matrix multiplexer JE2BEG3 MUX-16
assign JE2BEG3_input = {W6END0,W2END4,SS4END3,S2END4,E6END0,E2END4,N4END0,N2END4,N1END2,o_6to27,o_6to26,o_6to25,o_6to24,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG3 (
    .A0(JE2BEG3_input[0]),
    .A1(JE2BEG3_input[1]),
    .A2(JE2BEG3_input[2]),
    .A3(JE2BEG3_input[3]),
    .A4(JE2BEG3_input[4]),
    .A5(JE2BEG3_input[5]),
    .A6(JE2BEG3_input[6]),
    .A7(JE2BEG3_input[7]),
    .A8(JE2BEG3_input[8]),
    .A9(JE2BEG3_input[9]),
    .A10(JE2BEG3_input[10]),
    .A11(JE2BEG3_input[11]),
    .A12(JE2BEG3_input[12]),
    .A13(JE2BEG3_input[13]),
    .A14(JE2BEG3_input[14]),
    .A15(JE2BEG3_input[15]),
    .S0(ConfigBits[268+0]),
    .S0N(ConfigBits_N[268+0]),
    .S1(ConfigBits[268+1]),
    .S1N(ConfigBits_N[268+1]),
    .S2(ConfigBits[268+2]),
    .S2N(ConfigBits_N[268+2]),
    .S3(ConfigBits[268+3]),
    .S3N(ConfigBits_N[268+3]),
    .X(JE2BEG3)
);

 //switch matrix multiplexer JE2BEG4 MUX-16
assign JE2BEG4_input = {W1END1,S2END5,S1END3,S1END1,EE4END3,E2END5,E1END1,N2END5,N1END1,o_6to27,o_6to26,o_6to25,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG4 (
    .A0(JE2BEG4_input[0]),
    .A1(JE2BEG4_input[1]),
    .A2(JE2BEG4_input[2]),
    .A3(JE2BEG4_input[3]),
    .A4(JE2BEG4_input[4]),
    .A5(JE2BEG4_input[5]),
    .A6(JE2BEG4_input[6]),
    .A7(JE2BEG4_input[7]),
    .A8(JE2BEG4_input[8]),
    .A9(JE2BEG4_input[9]),
    .A10(JE2BEG4_input[10]),
    .A11(JE2BEG4_input[11]),
    .A12(JE2BEG4_input[12]),
    .A13(JE2BEG4_input[13]),
    .A14(JE2BEG4_input[14]),
    .A15(JE2BEG4_input[15]),
    .S0(ConfigBits[272+0]),
    .S0N(ConfigBits_N[272+0]),
    .S1(ConfigBits[272+1]),
    .S1N(ConfigBits_N[272+1]),
    .S2(ConfigBits[272+2]),
    .S2N(ConfigBits_N[272+2]),
    .S3(ConfigBits[272+3]),
    .S3N(ConfigBits_N[272+3]),
    .X(JE2BEG4)
);

 //switch matrix multiplexer JE2BEG5 MUX-16
assign JE2BEG5_input = {W1END2,S2END6,S1END2,S1END0,EE4END2,E2END6,E1END2,N2END6,N1END2,o_6to27,o_6to26,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG5 (
    .A0(JE2BEG5_input[0]),
    .A1(JE2BEG5_input[1]),
    .A2(JE2BEG5_input[2]),
    .A3(JE2BEG5_input[3]),
    .A4(JE2BEG5_input[4]),
    .A5(JE2BEG5_input[5]),
    .A6(JE2BEG5_input[6]),
    .A7(JE2BEG5_input[7]),
    .A8(JE2BEG5_input[8]),
    .A9(JE2BEG5_input[9]),
    .A10(JE2BEG5_input[10]),
    .A11(JE2BEG5_input[11]),
    .A12(JE2BEG5_input[12]),
    .A13(JE2BEG5_input[13]),
    .A14(JE2BEG5_input[14]),
    .A15(JE2BEG5_input[15]),
    .S0(ConfigBits[276+0]),
    .S0N(ConfigBits_N[276+0]),
    .S1(ConfigBits[276+1]),
    .S1N(ConfigBits_N[276+1]),
    .S2(ConfigBits[276+2]),
    .S2N(ConfigBits_N[276+2]),
    .S3(ConfigBits[276+3]),
    .S3N(ConfigBits_N[276+3]),
    .X(JE2BEG5)
);

 //switch matrix multiplexer JE2BEG6 MUX-16
assign JE2BEG6_input = {W1END3,S2END7,S1END3,S1END1,EE4END1,E2END7,E1END3,N2END7,N1END3,o_6to27,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG6 (
    .A0(JE2BEG6_input[0]),
    .A1(JE2BEG6_input[1]),
    .A2(JE2BEG6_input[2]),
    .A3(JE2BEG6_input[3]),
    .A4(JE2BEG6_input[4]),
    .A5(JE2BEG6_input[5]),
    .A6(JE2BEG6_input[6]),
    .A7(JE2BEG6_input[7]),
    .A8(JE2BEG6_input[8]),
    .A9(JE2BEG6_input[9]),
    .A10(JE2BEG6_input[10]),
    .A11(JE2BEG6_input[11]),
    .A12(JE2BEG6_input[12]),
    .A13(JE2BEG6_input[13]),
    .A14(JE2BEG6_input[14]),
    .A15(JE2BEG6_input[15]),
    .S0(ConfigBits[280+0]),
    .S0N(ConfigBits_N[280+0]),
    .S1(ConfigBits[280+1]),
    .S1N(ConfigBits_N[280+1]),
    .S2(ConfigBits[280+2]),
    .S2N(ConfigBits_N[280+2]),
    .S3(ConfigBits[280+3]),
    .S3N(ConfigBits_N[280+3]),
    .X(JE2BEG6)
);

 //switch matrix multiplexer JE2BEG7 MUX-16
assign JE2BEG7_input = {W1END0,S2END0,S1END2,S1END0,EE4END0,E2END0,E1END0,N2END0,N1END0,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JE2BEG7 (
    .A0(JE2BEG7_input[0]),
    .A1(JE2BEG7_input[1]),
    .A2(JE2BEG7_input[2]),
    .A3(JE2BEG7_input[3]),
    .A4(JE2BEG7_input[4]),
    .A5(JE2BEG7_input[5]),
    .A6(JE2BEG7_input[6]),
    .A7(JE2BEG7_input[7]),
    .A8(JE2BEG7_input[8]),
    .A9(JE2BEG7_input[9]),
    .A10(JE2BEG7_input[10]),
    .A11(JE2BEG7_input[11]),
    .A12(JE2BEG7_input[12]),
    .A13(JE2BEG7_input[13]),
    .A14(JE2BEG7_input[14]),
    .A15(JE2BEG7_input[15]),
    .S0(ConfigBits[284+0]),
    .S0N(ConfigBits_N[284+0]),
    .S1(ConfigBits[284+1]),
    .S1N(ConfigBits_N[284+1]),
    .S2(ConfigBits[284+2]),
    .S2N(ConfigBits_N[284+2]),
    .S3(ConfigBits[284+3]),
    .S3N(ConfigBits_N[284+3]),
    .X(JE2BEG7)
);

 //switch matrix multiplexer JS2BEG0 MUX-16
assign JS2BEG0_input = {W6END1,WW4END0,W2END1,S4END1,S2END1,E6END1,E2END1,E1END3,N2END1,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG0 (
    .A0(JS2BEG0_input[0]),
    .A1(JS2BEG0_input[1]),
    .A2(JS2BEG0_input[2]),
    .A3(JS2BEG0_input[3]),
    .A4(JS2BEG0_input[4]),
    .A5(JS2BEG0_input[5]),
    .A6(JS2BEG0_input[6]),
    .A7(JS2BEG0_input[7]),
    .A8(JS2BEG0_input[8]),
    .A9(JS2BEG0_input[9]),
    .A10(JS2BEG0_input[10]),
    .A11(JS2BEG0_input[11]),
    .A12(JS2BEG0_input[12]),
    .A13(JS2BEG0_input[13]),
    .A14(JS2BEG0_input[14]),
    .A15(JS2BEG0_input[15]),
    .S0(ConfigBits[288+0]),
    .S0N(ConfigBits_N[288+0]),
    .S1(ConfigBits[288+1]),
    .S1N(ConfigBits_N[288+1]),
    .S2(ConfigBits[288+2]),
    .S2N(ConfigBits_N[288+2]),
    .S3(ConfigBits[288+3]),
    .S3N(ConfigBits_N[288+3]),
    .X(JS2BEG0)
);

 //switch matrix multiplexer JS2BEG1 MUX-16
assign JS2BEG1_input = {W6END0,WW4END1,W2END2,S4END2,S2END2,E6END0,E2END2,E1END0,N2END2,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG1 (
    .A0(JS2BEG1_input[0]),
    .A1(JS2BEG1_input[1]),
    .A2(JS2BEG1_input[2]),
    .A3(JS2BEG1_input[3]),
    .A4(JS2BEG1_input[4]),
    .A5(JS2BEG1_input[5]),
    .A6(JS2BEG1_input[6]),
    .A7(JS2BEG1_input[7]),
    .A8(JS2BEG1_input[8]),
    .A9(JS2BEG1_input[9]),
    .A10(JS2BEG1_input[10]),
    .A11(JS2BEG1_input[11]),
    .A12(JS2BEG1_input[12]),
    .A13(JS2BEG1_input[13]),
    .A14(JS2BEG1_input[14]),
    .A15(JS2BEG1_input[15]),
    .S0(ConfigBits[292+0]),
    .S0N(ConfigBits_N[292+0]),
    .S1(ConfigBits[292+1]),
    .S1N(ConfigBits_N[292+1]),
    .S2(ConfigBits[292+2]),
    .S2N(ConfigBits_N[292+2]),
    .S3(ConfigBits[292+3]),
    .S3N(ConfigBits_N[292+3]),
    .X(JS2BEG1)
);

 //switch matrix multiplexer JS2BEG2 MUX-16
assign JS2BEG2_input = {W6END1,W2END3,S4END3,S2END3,E6END1,EE4END2,E2END3,E1END1,N2END3,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG2 (
    .A0(JS2BEG2_input[0]),
    .A1(JS2BEG2_input[1]),
    .A2(JS2BEG2_input[2]),
    .A3(JS2BEG2_input[3]),
    .A4(JS2BEG2_input[4]),
    .A5(JS2BEG2_input[5]),
    .A6(JS2BEG2_input[6]),
    .A7(JS2BEG2_input[7]),
    .A8(JS2BEG2_input[8]),
    .A9(JS2BEG2_input[9]),
    .A10(JS2BEG2_input[10]),
    .A11(JS2BEG2_input[11]),
    .A12(JS2BEG2_input[12]),
    .A13(JS2BEG2_input[13]),
    .A14(JS2BEG2_input[14]),
    .A15(JS2BEG2_input[15]),
    .S0(ConfigBits[296+0]),
    .S0N(ConfigBits_N[296+0]),
    .S1(ConfigBits[296+1]),
    .S1N(ConfigBits_N[296+1]),
    .S2(ConfigBits[296+2]),
    .S2N(ConfigBits_N[296+2]),
    .S3(ConfigBits[296+3]),
    .S3N(ConfigBits_N[296+3]),
    .X(JS2BEG2)
);

 //switch matrix multiplexer JS2BEG3 MUX-16
assign JS2BEG3_input = {W6END0,W2END4,S4END0,S2END4,E6END0,EE4END3,E2END4,E1END2,N2END4,o_6to27,o_6to26,o_6to25,o_6to24,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG3 (
    .A0(JS2BEG3_input[0]),
    .A1(JS2BEG3_input[1]),
    .A2(JS2BEG3_input[2]),
    .A3(JS2BEG3_input[3]),
    .A4(JS2BEG3_input[4]),
    .A5(JS2BEG3_input[5]),
    .A6(JS2BEG3_input[6]),
    .A7(JS2BEG3_input[7]),
    .A8(JS2BEG3_input[8]),
    .A9(JS2BEG3_input[9]),
    .A10(JS2BEG3_input[10]),
    .A11(JS2BEG3_input[11]),
    .A12(JS2BEG3_input[12]),
    .A13(JS2BEG3_input[13]),
    .A14(JS2BEG3_input[14]),
    .A15(JS2BEG3_input[15]),
    .S0(ConfigBits[300+0]),
    .S0N(ConfigBits_N[300+0]),
    .S1(ConfigBits[300+1]),
    .S1N(ConfigBits_N[300+1]),
    .S2(ConfigBits[300+2]),
    .S2N(ConfigBits_N[300+2]),
    .S3(ConfigBits[300+3]),
    .S3N(ConfigBits_N[300+3]),
    .X(JS2BEG3)
);

 //switch matrix multiplexer JS2BEG4 MUX-16
assign JS2BEG4_input = {W1END3,W1END1,SS4END3,S2END5,S1END1,E2END5,E1END1,N2END5,N1END1,o_6to27,o_6to26,o_6to25,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG4 (
    .A0(JS2BEG4_input[0]),
    .A1(JS2BEG4_input[1]),
    .A2(JS2BEG4_input[2]),
    .A3(JS2BEG4_input[3]),
    .A4(JS2BEG4_input[4]),
    .A5(JS2BEG4_input[5]),
    .A6(JS2BEG4_input[6]),
    .A7(JS2BEG4_input[7]),
    .A8(JS2BEG4_input[8]),
    .A9(JS2BEG4_input[9]),
    .A10(JS2BEG4_input[10]),
    .A11(JS2BEG4_input[11]),
    .A12(JS2BEG4_input[12]),
    .A13(JS2BEG4_input[13]),
    .A14(JS2BEG4_input[14]),
    .A15(JS2BEG4_input[15]),
    .S0(ConfigBits[304+0]),
    .S0N(ConfigBits_N[304+0]),
    .S1(ConfigBits[304+1]),
    .S1N(ConfigBits_N[304+1]),
    .S2(ConfigBits[304+2]),
    .S2N(ConfigBits_N[304+2]),
    .S3(ConfigBits[304+3]),
    .S3N(ConfigBits_N[304+3]),
    .X(JS2BEG4)
);

 //switch matrix multiplexer JS2BEG5 MUX-16
assign JS2BEG5_input = {W1END2,W1END0,SS4END2,S2END6,S1END2,E2END6,E1END2,N2END6,N1END2,o_6to27,o_6to26,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG5 (
    .A0(JS2BEG5_input[0]),
    .A1(JS2BEG5_input[1]),
    .A2(JS2BEG5_input[2]),
    .A3(JS2BEG5_input[3]),
    .A4(JS2BEG5_input[4]),
    .A5(JS2BEG5_input[5]),
    .A6(JS2BEG5_input[6]),
    .A7(JS2BEG5_input[7]),
    .A8(JS2BEG5_input[8]),
    .A9(JS2BEG5_input[9]),
    .A10(JS2BEG5_input[10]),
    .A11(JS2BEG5_input[11]),
    .A12(JS2BEG5_input[12]),
    .A13(JS2BEG5_input[13]),
    .A14(JS2BEG5_input[14]),
    .A15(JS2BEG5_input[15]),
    .S0(ConfigBits[308+0]),
    .S0N(ConfigBits_N[308+0]),
    .S1(ConfigBits[308+1]),
    .S1N(ConfigBits_N[308+1]),
    .S2(ConfigBits[308+2]),
    .S2N(ConfigBits_N[308+2]),
    .S3(ConfigBits[308+3]),
    .S3N(ConfigBits_N[308+3]),
    .X(JS2BEG5)
);

 //switch matrix multiplexer JS2BEG6 MUX-16
assign JS2BEG6_input = {W1END3,W1END1,SS4END1,S2END7,S1END3,E2END7,E1END3,N2END7,N1END3,o_6to27,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG6 (
    .A0(JS2BEG6_input[0]),
    .A1(JS2BEG6_input[1]),
    .A2(JS2BEG6_input[2]),
    .A3(JS2BEG6_input[3]),
    .A4(JS2BEG6_input[4]),
    .A5(JS2BEG6_input[5]),
    .A6(JS2BEG6_input[6]),
    .A7(JS2BEG6_input[7]),
    .A8(JS2BEG6_input[8]),
    .A9(JS2BEG6_input[9]),
    .A10(JS2BEG6_input[10]),
    .A11(JS2BEG6_input[11]),
    .A12(JS2BEG6_input[12]),
    .A13(JS2BEG6_input[13]),
    .A14(JS2BEG6_input[14]),
    .A15(JS2BEG6_input[15]),
    .S0(ConfigBits[312+0]),
    .S0N(ConfigBits_N[312+0]),
    .S1(ConfigBits[312+1]),
    .S1N(ConfigBits_N[312+1]),
    .S2(ConfigBits[312+2]),
    .S2N(ConfigBits_N[312+2]),
    .S3(ConfigBits[312+3]),
    .S3N(ConfigBits_N[312+3]),
    .X(JS2BEG6)
);

 //switch matrix multiplexer JS2BEG7 MUX-16
assign JS2BEG7_input = {W1END2,W1END0,SS4END0,S2END0,S1END0,E2END0,E1END0,N2END0,N1END0,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JS2BEG7 (
    .A0(JS2BEG7_input[0]),
    .A1(JS2BEG7_input[1]),
    .A2(JS2BEG7_input[2]),
    .A3(JS2BEG7_input[3]),
    .A4(JS2BEG7_input[4]),
    .A5(JS2BEG7_input[5]),
    .A6(JS2BEG7_input[6]),
    .A7(JS2BEG7_input[7]),
    .A8(JS2BEG7_input[8]),
    .A9(JS2BEG7_input[9]),
    .A10(JS2BEG7_input[10]),
    .A11(JS2BEG7_input[11]),
    .A12(JS2BEG7_input[12]),
    .A13(JS2BEG7_input[13]),
    .A14(JS2BEG7_input[14]),
    .A15(JS2BEG7_input[15]),
    .S0(ConfigBits[316+0]),
    .S0N(ConfigBits_N[316+0]),
    .S1(ConfigBits[316+1]),
    .S1N(ConfigBits_N[316+1]),
    .S2(ConfigBits[316+2]),
    .S2N(ConfigBits_N[316+2]),
    .S3(ConfigBits[316+3]),
    .S3N(ConfigBits_N[316+3]),
    .X(JS2BEG7)
);

 //switch matrix multiplexer JW2BEG0 MUX-16
assign JW2BEG0_input = {W6END1,W2END1,SS4END0,S4END1,S2END1,E6END1,E2END1,N2END1,N1END3,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG0 (
    .A0(JW2BEG0_input[0]),
    .A1(JW2BEG0_input[1]),
    .A2(JW2BEG0_input[2]),
    .A3(JW2BEG0_input[3]),
    .A4(JW2BEG0_input[4]),
    .A5(JW2BEG0_input[5]),
    .A6(JW2BEG0_input[6]),
    .A7(JW2BEG0_input[7]),
    .A8(JW2BEG0_input[8]),
    .A9(JW2BEG0_input[9]),
    .A10(JW2BEG0_input[10]),
    .A11(JW2BEG0_input[11]),
    .A12(JW2BEG0_input[12]),
    .A13(JW2BEG0_input[13]),
    .A14(JW2BEG0_input[14]),
    .A15(JW2BEG0_input[15]),
    .S0(ConfigBits[320+0]),
    .S0N(ConfigBits_N[320+0]),
    .S1(ConfigBits[320+1]),
    .S1N(ConfigBits_N[320+1]),
    .S2(ConfigBits[320+2]),
    .S2N(ConfigBits_N[320+2]),
    .S3(ConfigBits[320+3]),
    .S3N(ConfigBits_N[320+3]),
    .X(JW2BEG0)
);

 //switch matrix multiplexer JW2BEG1 MUX-16
assign JW2BEG1_input = {W6END0,W2END2,SS4END1,S4END2,S2END2,E6END0,E2END2,N2END2,N1END0,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG1 (
    .A0(JW2BEG1_input[0]),
    .A1(JW2BEG1_input[1]),
    .A2(JW2BEG1_input[2]),
    .A3(JW2BEG1_input[3]),
    .A4(JW2BEG1_input[4]),
    .A5(JW2BEG1_input[5]),
    .A6(JW2BEG1_input[6]),
    .A7(JW2BEG1_input[7]),
    .A8(JW2BEG1_input[8]),
    .A9(JW2BEG1_input[9]),
    .A10(JW2BEG1_input[10]),
    .A11(JW2BEG1_input[11]),
    .A12(JW2BEG1_input[12]),
    .A13(JW2BEG1_input[13]),
    .A14(JW2BEG1_input[14]),
    .A15(JW2BEG1_input[15]),
    .S0(ConfigBits[324+0]),
    .S0N(ConfigBits_N[324+0]),
    .S1(ConfigBits[324+1]),
    .S1N(ConfigBits_N[324+1]),
    .S2(ConfigBits[324+2]),
    .S2N(ConfigBits_N[324+2]),
    .S3(ConfigBits[324+3]),
    .S3N(ConfigBits_N[324+3]),
    .X(JW2BEG1)
);

 //switch matrix multiplexer JW2BEG2 MUX-16
assign JW2BEG2_input = {W6END1,W2END3,S4END3,S2END3,E6END1,E2END3,NN4END2,N2END3,N1END1,o_6to27,o_6to26,o_6to25,o_6to24,o_6to23,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG2 (
    .A0(JW2BEG2_input[0]),
    .A1(JW2BEG2_input[1]),
    .A2(JW2BEG2_input[2]),
    .A3(JW2BEG2_input[3]),
    .A4(JW2BEG2_input[4]),
    .A5(JW2BEG2_input[5]),
    .A6(JW2BEG2_input[6]),
    .A7(JW2BEG2_input[7]),
    .A8(JW2BEG2_input[8]),
    .A9(JW2BEG2_input[9]),
    .A10(JW2BEG2_input[10]),
    .A11(JW2BEG2_input[11]),
    .A12(JW2BEG2_input[12]),
    .A13(JW2BEG2_input[13]),
    .A14(JW2BEG2_input[14]),
    .A15(JW2BEG2_input[15]),
    .S0(ConfigBits[328+0]),
    .S0N(ConfigBits_N[328+0]),
    .S1(ConfigBits[328+1]),
    .S1N(ConfigBits_N[328+1]),
    .S2(ConfigBits[328+2]),
    .S2N(ConfigBits_N[328+2]),
    .S3(ConfigBits[328+3]),
    .S3N(ConfigBits_N[328+3]),
    .X(JW2BEG2)
);

 //switch matrix multiplexer JW2BEG3 MUX-16
assign JW2BEG3_input = {W6END0,W2END4,S4END0,S2END4,E6END0,E2END4,NN4END3,N2END4,N1END2,o_6to27,o_6to26,o_6to25,o_6to24,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG3 (
    .A0(JW2BEG3_input[0]),
    .A1(JW2BEG3_input[1]),
    .A2(JW2BEG3_input[2]),
    .A3(JW2BEG3_input[3]),
    .A4(JW2BEG3_input[4]),
    .A5(JW2BEG3_input[5]),
    .A6(JW2BEG3_input[6]),
    .A7(JW2BEG3_input[7]),
    .A8(JW2BEG3_input[8]),
    .A9(JW2BEG3_input[9]),
    .A10(JW2BEG3_input[10]),
    .A11(JW2BEG3_input[11]),
    .A12(JW2BEG3_input[12]),
    .A13(JW2BEG3_input[13]),
    .A14(JW2BEG3_input[14]),
    .A15(JW2BEG3_input[15]),
    .S0(ConfigBits[332+0]),
    .S0N(ConfigBits_N[332+0]),
    .S1(ConfigBits[332+1]),
    .S1N(ConfigBits_N[332+1]),
    .S2(ConfigBits[332+2]),
    .S2N(ConfigBits_N[332+2]),
    .S3(ConfigBits[332+3]),
    .S3N(ConfigBits_N[332+3]),
    .X(JW2BEG3)
);

 //switch matrix multiplexer JW2BEG4 MUX-16
assign JW2BEG4_input = {WW4END3,W1END1,S2END5,S1END3,S1END1,E2END5,E1END1,N2END5,N1END1,o_6to27,o_6to26,o_6to25,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG4 (
    .A0(JW2BEG4_input[0]),
    .A1(JW2BEG4_input[1]),
    .A2(JW2BEG4_input[2]),
    .A3(JW2BEG4_input[3]),
    .A4(JW2BEG4_input[4]),
    .A5(JW2BEG4_input[5]),
    .A6(JW2BEG4_input[6]),
    .A7(JW2BEG4_input[7]),
    .A8(JW2BEG4_input[8]),
    .A9(JW2BEG4_input[9]),
    .A10(JW2BEG4_input[10]),
    .A11(JW2BEG4_input[11]),
    .A12(JW2BEG4_input[12]),
    .A13(JW2BEG4_input[13]),
    .A14(JW2BEG4_input[14]),
    .A15(JW2BEG4_input[15]),
    .S0(ConfigBits[336+0]),
    .S0N(ConfigBits_N[336+0]),
    .S1(ConfigBits[336+1]),
    .S1N(ConfigBits_N[336+1]),
    .S2(ConfigBits[336+2]),
    .S2N(ConfigBits_N[336+2]),
    .S3(ConfigBits[336+3]),
    .S3N(ConfigBits_N[336+3]),
    .X(JW2BEG4)
);

 //switch matrix multiplexer JW2BEG5 MUX-16
assign JW2BEG5_input = {WW4END2,W1END2,S2END6,S1END2,S1END0,E2END6,E1END2,N2END6,N1END2,o_6to27,o_6to26,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG5 (
    .A0(JW2BEG5_input[0]),
    .A1(JW2BEG5_input[1]),
    .A2(JW2BEG5_input[2]),
    .A3(JW2BEG5_input[3]),
    .A4(JW2BEG5_input[4]),
    .A5(JW2BEG5_input[5]),
    .A6(JW2BEG5_input[6]),
    .A7(JW2BEG5_input[7]),
    .A8(JW2BEG5_input[8]),
    .A9(JW2BEG5_input[9]),
    .A10(JW2BEG5_input[10]),
    .A11(JW2BEG5_input[11]),
    .A12(JW2BEG5_input[12]),
    .A13(JW2BEG5_input[13]),
    .A14(JW2BEG5_input[14]),
    .A15(JW2BEG5_input[15]),
    .S0(ConfigBits[340+0]),
    .S0N(ConfigBits_N[340+0]),
    .S1(ConfigBits[340+1]),
    .S1N(ConfigBits_N[340+1]),
    .S2(ConfigBits[340+2]),
    .S2N(ConfigBits_N[340+2]),
    .S3(ConfigBits[340+3]),
    .S3N(ConfigBits_N[340+3]),
    .X(JW2BEG5)
);

 //switch matrix multiplexer JW2BEG6 MUX-16
assign JW2BEG6_input = {WW4END1,W1END3,S2END7,S1END3,S1END1,E2END7,E1END3,N2END7,N1END3,o_6to27,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG6 (
    .A0(JW2BEG6_input[0]),
    .A1(JW2BEG6_input[1]),
    .A2(JW2BEG6_input[2]),
    .A3(JW2BEG6_input[3]),
    .A4(JW2BEG6_input[4]),
    .A5(JW2BEG6_input[5]),
    .A6(JW2BEG6_input[6]),
    .A7(JW2BEG6_input[7]),
    .A8(JW2BEG6_input[8]),
    .A9(JW2BEG6_input[9]),
    .A10(JW2BEG6_input[10]),
    .A11(JW2BEG6_input[11]),
    .A12(JW2BEG6_input[12]),
    .A13(JW2BEG6_input[13]),
    .A14(JW2BEG6_input[14]),
    .A15(JW2BEG6_input[15]),
    .S0(ConfigBits[344+0]),
    .S0N(ConfigBits_N[344+0]),
    .S1(ConfigBits[344+1]),
    .S1N(ConfigBits_N[344+1]),
    .S2(ConfigBits[344+2]),
    .S2N(ConfigBits_N[344+2]),
    .S3(ConfigBits[344+3]),
    .S3N(ConfigBits_N[344+3]),
    .X(JW2BEG6)
);

 //switch matrix multiplexer JW2BEG7 MUX-16
assign JW2BEG7_input = {WW4END0,W1END0,S2END0,S1END2,S1END0,E2END0,E1END0,N2END0,N1END0,o_6to26,o_6to25,o_6to24,o_6to23,o_6to22,o_6to21,o_6to20};
cus_mux161_buf inst_cus_mux161_buf_JW2BEG7 (
    .A0(JW2BEG7_input[0]),
    .A1(JW2BEG7_input[1]),
    .A2(JW2BEG7_input[2]),
    .A3(JW2BEG7_input[3]),
    .A4(JW2BEG7_input[4]),
    .A5(JW2BEG7_input[5]),
    .A6(JW2BEG7_input[6]),
    .A7(JW2BEG7_input[7]),
    .A8(JW2BEG7_input[8]),
    .A9(JW2BEG7_input[9]),
    .A10(JW2BEG7_input[10]),
    .A11(JW2BEG7_input[11]),
    .A12(JW2BEG7_input[12]),
    .A13(JW2BEG7_input[13]),
    .A14(JW2BEG7_input[14]),
    .A15(JW2BEG7_input[15]),
    .S0(ConfigBits[348+0]),
    .S0N(ConfigBits_N[348+0]),
    .S1(ConfigBits[348+1]),
    .S1N(ConfigBits_N[348+1]),
    .S2(ConfigBits[348+2]),
    .S2N(ConfigBits_N[348+2]),
    .S3(ConfigBits[348+3]),
    .S3N(ConfigBits_N[348+3]),
    .X(JW2BEG7)
);

 //switch matrix multiplexer J_l_AB_BEG0 MUX-4
assign J_l_AB_BEG0_input = {JN2END1,WW4END0,S4END3,NN4END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG0 (
    .A0(J_l_AB_BEG0_input[0]),
    .A1(J_l_AB_BEG0_input[1]),
    .A2(J_l_AB_BEG0_input[2]),
    .A3(J_l_AB_BEG0_input[3]),
    .S0(ConfigBits[352+0]),
    .S0N(ConfigBits_N[352+0]),
    .S1(ConfigBits[352+1]),
    .S1N(ConfigBits_N[352+1]),
    .X(J_l_AB_BEG0)
);

 //switch matrix multiplexer J_l_AB_BEG1 MUX-4
assign J_l_AB_BEG1_input = {JE2END1,W2END7,S4END2,EE4END2};
cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG1 (
    .A0(J_l_AB_BEG1_input[0]),
    .A1(J_l_AB_BEG1_input[1]),
    .A2(J_l_AB_BEG1_input[2]),
    .A3(J_l_AB_BEG1_input[3]),
    .S0(ConfigBits[354+0]),
    .S0N(ConfigBits_N[354+0]),
    .S1(ConfigBits[354+1]),
    .S1N(ConfigBits_N[354+1]),
    .X(J_l_AB_BEG1)
);

 //switch matrix multiplexer J_l_AB_BEG2 MUX-4
assign J_l_AB_BEG2_input = {JS2END1,W6END1,E6END1,N4END1};
cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG2 (
    .A0(J_l_AB_BEG2_input[0]),
    .A1(J_l_AB_BEG2_input[1]),
    .A2(J_l_AB_BEG2_input[2]),
    .A3(J_l_AB_BEG2_input[3]),
    .S0(ConfigBits[356+0]),
    .S0N(ConfigBits_N[356+0]),
    .S1(ConfigBits[356+1]),
    .S1N(ConfigBits_N[356+1]),
    .X(J_l_AB_BEG2)
);

 //switch matrix multiplexer J_l_AB_BEG3 MUX-4
assign J_l_AB_BEG3_input = {JW2END1,S4END0,E6END0,N4END0};
cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG3 (
    .A0(J_l_AB_BEG3_input[0]),
    .A1(J_l_AB_BEG3_input[1]),
    .A2(J_l_AB_BEG3_input[2]),
    .A3(J_l_AB_BEG3_input[3]),
    .S0(ConfigBits[358+0]),
    .S0N(ConfigBits_N[358+0]),
    .S1(ConfigBits[358+1]),
    .S1N(ConfigBits_N[358+1]),
    .X(J_l_AB_BEG3)
);

 //switch matrix multiplexer J_l_CD_BEG0 MUX-4
assign J_l_CD_BEG0_input = {JN2END2,WW4END2,SS4END3,E2END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG0 (
    .A0(J_l_CD_BEG0_input[0]),
    .A1(J_l_CD_BEG0_input[1]),
    .A2(J_l_CD_BEG0_input[2]),
    .A3(J_l_CD_BEG0_input[3]),
    .S0(ConfigBits[360+0]),
    .S0N(ConfigBits_N[360+0]),
    .S1(ConfigBits[360+1]),
    .S1N(ConfigBits_N[360+1]),
    .X(J_l_CD_BEG0)
);

 //switch matrix multiplexer J_l_CD_BEG1 MUX-4
assign J_l_CD_BEG1_input = {JE2END2,W2END7,E2END2,N4END2};
cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG1 (
    .A0(J_l_CD_BEG1_input[0]),
    .A1(J_l_CD_BEG1_input[1]),
    .A2(J_l_CD_BEG1_input[2]),
    .A3(J_l_CD_BEG1_input[3]),
    .S0(ConfigBits[362+0]),
    .S0N(ConfigBits_N[362+0]),
    .S1(ConfigBits[362+1]),
    .S1N(ConfigBits_N[362+1]),
    .X(J_l_CD_BEG1)
);

 //switch matrix multiplexer J_l_CD_BEG2 MUX-4
assign J_l_CD_BEG2_input = {JS2END2,S4END1,EE4END1,NN4END1};
cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG2 (
    .A0(J_l_CD_BEG2_input[0]),
    .A1(J_l_CD_BEG2_input[1]),
    .A2(J_l_CD_BEG2_input[2]),
    .A3(J_l_CD_BEG2_input[3]),
    .S0(ConfigBits[364+0]),
    .S0N(ConfigBits_N[364+0]),
    .S1(ConfigBits[364+1]),
    .S1N(ConfigBits_N[364+1]),
    .X(J_l_CD_BEG2)
);

 //switch matrix multiplexer J_l_CD_BEG3 MUX-4
assign J_l_CD_BEG3_input = {JW2END2,W6END0,SS4END0,N4END0};
cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG3 (
    .A0(J_l_CD_BEG3_input[0]),
    .A1(J_l_CD_BEG3_input[1]),
    .A2(J_l_CD_BEG3_input[2]),
    .A3(J_l_CD_BEG3_input[3]),
    .S0(ConfigBits[366+0]),
    .S0N(ConfigBits_N[366+0]),
    .S1(ConfigBits[366+1]),
    .S1N(ConfigBits_N[366+1]),
    .X(J_l_CD_BEG3)
);

 //switch matrix multiplexer J_l_EF_BEG0 MUX-4
assign J_l_EF_BEG0_input = {JN2END3,W2END3,E2END3,N4END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG0 (
    .A0(J_l_EF_BEG0_input[0]),
    .A1(J_l_EF_BEG0_input[1]),
    .A2(J_l_EF_BEG0_input[2]),
    .A3(J_l_EF_BEG0_input[3]),
    .S0(ConfigBits[368+0]),
    .S0N(ConfigBits_N[368+0]),
    .S1(ConfigBits[368+1]),
    .S1N(ConfigBits_N[368+1]),
    .X(J_l_EF_BEG0)
);

 //switch matrix multiplexer J_l_EF_BEG1 MUX-4
assign J_l_EF_BEG1_input = {JE2END3,S4END2,E2END2,NN4END2};
cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG1 (
    .A0(J_l_EF_BEG1_input[0]),
    .A1(J_l_EF_BEG1_input[1]),
    .A2(J_l_EF_BEG1_input[2]),
    .A3(J_l_EF_BEG1_input[3]),
    .S0(ConfigBits[370+0]),
    .S0N(ConfigBits_N[370+0]),
    .S1(ConfigBits[370+1]),
    .S1N(ConfigBits_N[370+1]),
    .X(J_l_EF_BEG1)
);

 //switch matrix multiplexer J_l_EF_BEG2 MUX-4
assign J_l_EF_BEG2_input = {JS2END3,W2END4,SS4END1,N4END1};
cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG2 (
    .A0(J_l_EF_BEG2_input[0]),
    .A1(J_l_EF_BEG2_input[1]),
    .A2(J_l_EF_BEG2_input[2]),
    .A3(J_l_EF_BEG2_input[3]),
    .S0(ConfigBits[372+0]),
    .S0N(ConfigBits_N[372+0]),
    .S1(ConfigBits[372+1]),
    .S1N(ConfigBits_N[372+1]),
    .X(J_l_EF_BEG2)
);

 //switch matrix multiplexer J_l_EF_BEG3 MUX-4
assign J_l_EF_BEG3_input = {JW2END3,WW4END1,S4END0,EE4END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG3 (
    .A0(J_l_EF_BEG3_input[0]),
    .A1(J_l_EF_BEG3_input[1]),
    .A2(J_l_EF_BEG3_input[2]),
    .A3(J_l_EF_BEG3_input[3]),
    .S0(ConfigBits[374+0]),
    .S0N(ConfigBits_N[374+0]),
    .S1(ConfigBits[374+1]),
    .S1N(ConfigBits_N[374+1]),
    .X(J_l_EF_BEG3)
);

 //switch matrix multiplexer J_l_GH_BEG0 MUX-4
assign J_l_GH_BEG0_input = {JN2END4,S4END3,EE4END0,N4END3};
cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG0 (
    .A0(J_l_GH_BEG0_input[0]),
    .A1(J_l_GH_BEG0_input[1]),
    .A2(J_l_GH_BEG0_input[2]),
    .A3(J_l_GH_BEG0_input[3]),
    .S0(ConfigBits[376+0]),
    .S0N(ConfigBits_N[376+0]),
    .S1(ConfigBits[376+1]),
    .S1N(ConfigBits_N[376+1]),
    .X(J_l_GH_BEG0)
);

 //switch matrix multiplexer J_l_GH_BEG1 MUX-4
assign J_l_GH_BEG1_input = {JE2END4,W2END2,SS4END2,N4END2};
cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG1 (
    .A0(J_l_GH_BEG1_input[0]),
    .A1(J_l_GH_BEG1_input[1]),
    .A2(J_l_GH_BEG1_input[2]),
    .A3(J_l_GH_BEG1_input[3]),
    .S0(ConfigBits[378+0]),
    .S0N(ConfigBits_N[378+0]),
    .S1(ConfigBits[378+1]),
    .S1N(ConfigBits_N[378+1]),
    .X(J_l_GH_BEG1)
);

 //switch matrix multiplexer J_l_GH_BEG2 MUX-4
assign J_l_GH_BEG2_input = {JS2END4,WW4END3,S4END1,E6END1};
cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG2 (
    .A0(J_l_GH_BEG2_input[0]),
    .A1(J_l_GH_BEG2_input[1]),
    .A2(J_l_GH_BEG2_input[2]),
    .A3(J_l_GH_BEG2_input[3]),
    .S0(ConfigBits[380+0]),
    .S0N(ConfigBits_N[380+0]),
    .S1(ConfigBits[380+1]),
    .S1N(ConfigBits_N[380+1]),
    .X(J_l_GH_BEG2)
);

 //switch matrix multiplexer J_l_GH_BEG3 MUX-4
assign J_l_GH_BEG3_input = {JW2END4,W2END0,E6END0,NN4END0};
cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG3 (
    .A0(J_l_GH_BEG3_input[0]),
    .A1(J_l_GH_BEG3_input[1]),
    .A2(J_l_GH_BEG3_input[2]),
    .A3(J_l_GH_BEG3_input[3]),
    .S0(ConfigBits[382+0]),
    .S0N(ConfigBits_N[382+0]),
    .S1(ConfigBits[382+1]),
    .S1N(ConfigBits_N[382+1]),
    .X(J_l_GH_BEG3)
);


assign DEBUG_select_i_2to60         = ConfigBits[1:0];
assign DEBUG_select_i_2to61         = ConfigBits[3:2];
assign DEBUG_select_i_2to62         = ConfigBits[5:4];
assign DEBUG_select_i_2to63         = ConfigBits[7:6];
assign DEBUG_select_i_2to64         = ConfigBits[9:8];
assign DEBUG_select_i_2to65         = ConfigBits[11:10];
assign DEBUG_select_i_2to66         = ConfigBits[13:12];
assign DEBUG_select_i_2to67         = ConfigBits[15:14];
assign DEBUG_select_N1BEG0          = ConfigBits[17:16];
assign DEBUG_select_N1BEG1          = ConfigBits[19:18];
assign DEBUG_select_N1BEG2          = ConfigBits[21:20];
assign DEBUG_select_N1BEG3          = ConfigBits[23:22];
assign DEBUG_select_N4BEG0          = ConfigBits[25:24];
assign DEBUG_select_N4BEG1          = ConfigBits[27:26];
assign DEBUG_select_N4BEG2          = ConfigBits[29:28];
assign DEBUG_select_N4BEG3          = ConfigBits[31:30];
assign DEBUG_select_NN4BEG0         = ConfigBits[34:32];
assign DEBUG_select_NN4BEG1         = ConfigBits[37:35];
assign DEBUG_select_NN4BEG2         = ConfigBits[40:38];
assign DEBUG_select_NN4BEG3         = ConfigBits[43:41];
assign DEBUG_select_E1BEG0          = ConfigBits[45:44];
assign DEBUG_select_E1BEG1          = ConfigBits[47:46];
assign DEBUG_select_E1BEG2          = ConfigBits[49:48];
assign DEBUG_select_E1BEG3          = ConfigBits[51:50];
assign DEBUG_select_EE4BEG0         = ConfigBits[54:52];
assign DEBUG_select_EE4BEG1         = ConfigBits[57:55];
assign DEBUG_select_EE4BEG2         = ConfigBits[60:58];
assign DEBUG_select_EE4BEG3         = ConfigBits[63:61];
assign DEBUG_select_E6BEG0          = ConfigBits[67:64];
assign DEBUG_select_E6BEG1          = ConfigBits[71:68];
assign DEBUG_select_S1BEG0          = ConfigBits[73:72];
assign DEBUG_select_S1BEG1          = ConfigBits[75:74];
assign DEBUG_select_S1BEG2          = ConfigBits[77:76];
assign DEBUG_select_S1BEG3          = ConfigBits[79:78];
assign DEBUG_select_S4BEG0          = ConfigBits[81:80];
assign DEBUG_select_S4BEG1          = ConfigBits[83:82];
assign DEBUG_select_S4BEG2          = ConfigBits[85:84];
assign DEBUG_select_S4BEG3          = ConfigBits[87:86];
assign DEBUG_select_SS4BEG0         = ConfigBits[90:88];
assign DEBUG_select_SS4BEG1         = ConfigBits[93:91];
assign DEBUG_select_SS4BEG2         = ConfigBits[96:94];
assign DEBUG_select_SS4BEG3         = ConfigBits[99:97];
assign DEBUG_select_W1BEG0          = ConfigBits[101:100];
assign DEBUG_select_W1BEG1          = ConfigBits[103:102];
assign DEBUG_select_W1BEG2          = ConfigBits[105:104];
assign DEBUG_select_W1BEG3          = ConfigBits[107:106];
assign DEBUG_select_WW4BEG0         = ConfigBits[110:108];
assign DEBUG_select_WW4BEG1         = ConfigBits[113:111];
assign DEBUG_select_WW4BEG2         = ConfigBits[116:114];
assign DEBUG_select_WW4BEG3         = ConfigBits[119:117];
assign DEBUG_select_W6BEG0          = ConfigBits[123:120];
assign DEBUG_select_W6BEG1          = ConfigBits[127:124];
assign DEBUG_select_J2MID_ABa_BEG0  = ConfigBits[129:128];
assign DEBUG_select_J2MID_ABa_BEG1  = ConfigBits[131:130];
assign DEBUG_select_J2MID_ABa_BEG2  = ConfigBits[133:132];
assign DEBUG_select_J2MID_ABa_BEG3  = ConfigBits[135:134];
assign DEBUG_select_J2MID_CDa_BEG0  = ConfigBits[137:136];
assign DEBUG_select_J2MID_CDa_BEG1  = ConfigBits[139:138];
assign DEBUG_select_J2MID_CDa_BEG2  = ConfigBits[141:140];
assign DEBUG_select_J2MID_CDa_BEG3  = ConfigBits[143:142];
assign DEBUG_select_J2MID_EFa_BEG0  = ConfigBits[145:144];
assign DEBUG_select_J2MID_EFa_BEG1  = ConfigBits[147:146];
assign DEBUG_select_J2MID_EFa_BEG2  = ConfigBits[149:148];
assign DEBUG_select_J2MID_EFa_BEG3  = ConfigBits[151:150];
assign DEBUG_select_J2MID_GHa_BEG0  = ConfigBits[153:152];
assign DEBUG_select_J2MID_GHa_BEG1  = ConfigBits[155:154];
assign DEBUG_select_J2MID_GHa_BEG2  = ConfigBits[157:156];
assign DEBUG_select_J2MID_GHa_BEG3  = ConfigBits[159:158];
assign DEBUG_select_J2MID_ABb_BEG0  = ConfigBits[161:160];
assign DEBUG_select_J2MID_ABb_BEG1  = ConfigBits[163:162];
assign DEBUG_select_J2MID_ABb_BEG2  = ConfigBits[165:164];
assign DEBUG_select_J2MID_ABb_BEG3  = ConfigBits[167:166];
assign DEBUG_select_J2MID_CDb_BEG0  = ConfigBits[169:168];
assign DEBUG_select_J2MID_CDb_BEG1  = ConfigBits[171:170];
assign DEBUG_select_J2MID_CDb_BEG2  = ConfigBits[173:172];
assign DEBUG_select_J2MID_CDb_BEG3  = ConfigBits[175:174];
assign DEBUG_select_J2MID_EFb_BEG0  = ConfigBits[177:176];
assign DEBUG_select_J2MID_EFb_BEG1  = ConfigBits[179:178];
assign DEBUG_select_J2MID_EFb_BEG2  = ConfigBits[181:180];
assign DEBUG_select_J2MID_EFb_BEG3  = ConfigBits[183:182];
assign DEBUG_select_J2MID_GHb_BEG0  = ConfigBits[185:184];
assign DEBUG_select_J2MID_GHb_BEG1  = ConfigBits[187:186];
assign DEBUG_select_J2MID_GHb_BEG2  = ConfigBits[189:188];
assign DEBUG_select_J2MID_GHb_BEG3  = ConfigBits[191:190];
assign DEBUG_select_J2END_AB_BEG0   = ConfigBits[193:192];
assign DEBUG_select_J2END_AB_BEG1   = ConfigBits[195:194];
assign DEBUG_select_J2END_AB_BEG2   = ConfigBits[197:196];
assign DEBUG_select_J2END_AB_BEG3   = ConfigBits[199:198];
assign DEBUG_select_J2END_CD_BEG0   = ConfigBits[201:200];
assign DEBUG_select_J2END_CD_BEG1   = ConfigBits[203:202];
assign DEBUG_select_J2END_CD_BEG2   = ConfigBits[205:204];
assign DEBUG_select_J2END_CD_BEG3   = ConfigBits[207:206];
assign DEBUG_select_J2END_EF_BEG0   = ConfigBits[209:208];
assign DEBUG_select_J2END_EF_BEG1   = ConfigBits[211:210];
assign DEBUG_select_J2END_EF_BEG2   = ConfigBits[213:212];
assign DEBUG_select_J2END_EF_BEG3   = ConfigBits[215:214];
assign DEBUG_select_J2END_GH_BEG0   = ConfigBits[217:216];
assign DEBUG_select_J2END_GH_BEG1   = ConfigBits[219:218];
assign DEBUG_select_J2END_GH_BEG2   = ConfigBits[221:220];
assign DEBUG_select_J2END_GH_BEG3   = ConfigBits[223:222];
assign DEBUG_select_JN2BEG0         = ConfigBits[227:224];
assign DEBUG_select_JN2BEG1         = ConfigBits[231:228];
assign DEBUG_select_JN2BEG2         = ConfigBits[235:232];
assign DEBUG_select_JN2BEG3         = ConfigBits[239:236];
assign DEBUG_select_JN2BEG4         = ConfigBits[243:240];
assign DEBUG_select_JN2BEG5         = ConfigBits[247:244];
assign DEBUG_select_JN2BEG6         = ConfigBits[251:248];
assign DEBUG_select_JN2BEG7         = ConfigBits[255:252];
assign DEBUG_select_JE2BEG0         = ConfigBits[259:256];
assign DEBUG_select_JE2BEG1         = ConfigBits[263:260];
assign DEBUG_select_JE2BEG2         = ConfigBits[267:264];
assign DEBUG_select_JE2BEG3         = ConfigBits[271:268];
assign DEBUG_select_JE2BEG4         = ConfigBits[275:272];
assign DEBUG_select_JE2BEG5         = ConfigBits[279:276];
assign DEBUG_select_JE2BEG6         = ConfigBits[283:280];
assign DEBUG_select_JE2BEG7         = ConfigBits[287:284];
assign DEBUG_select_JS2BEG0         = ConfigBits[291:288];
assign DEBUG_select_JS2BEG1         = ConfigBits[295:292];
assign DEBUG_select_JS2BEG2         = ConfigBits[299:296];
assign DEBUG_select_JS2BEG3         = ConfigBits[303:300];
assign DEBUG_select_JS2BEG4         = ConfigBits[307:304];
assign DEBUG_select_JS2BEG5         = ConfigBits[311:308];
assign DEBUG_select_JS2BEG6         = ConfigBits[315:312];
assign DEBUG_select_JS2BEG7         = ConfigBits[319:316];
assign DEBUG_select_JW2BEG0         = ConfigBits[323:320];
assign DEBUG_select_JW2BEG1         = ConfigBits[327:324];
assign DEBUG_select_JW2BEG2         = ConfigBits[331:328];
assign DEBUG_select_JW2BEG3         = ConfigBits[335:332];
assign DEBUG_select_JW2BEG4         = ConfigBits[339:336];
assign DEBUG_select_JW2BEG5         = ConfigBits[343:340];
assign DEBUG_select_JW2BEG6         = ConfigBits[347:344];
assign DEBUG_select_JW2BEG7         = ConfigBits[351:348];
assign DEBUG_select_J_l_AB_BEG0     = ConfigBits[353:352];
assign DEBUG_select_J_l_AB_BEG1     = ConfigBits[355:354];
assign DEBUG_select_J_l_AB_BEG2     = ConfigBits[357:356];
assign DEBUG_select_J_l_AB_BEG3     = ConfigBits[359:358];
assign DEBUG_select_J_l_CD_BEG0     = ConfigBits[361:360];
assign DEBUG_select_J_l_CD_BEG1     = ConfigBits[363:362];
assign DEBUG_select_J_l_CD_BEG2     = ConfigBits[365:364];
assign DEBUG_select_J_l_CD_BEG3     = ConfigBits[367:366];
assign DEBUG_select_J_l_EF_BEG0     = ConfigBits[369:368];
assign DEBUG_select_J_l_EF_BEG1     = ConfigBits[371:370];
assign DEBUG_select_J_l_EF_BEG2     = ConfigBits[373:372];
assign DEBUG_select_J_l_EF_BEG3     = ConfigBits[375:374];
assign DEBUG_select_J_l_GH_BEG0     = ConfigBits[377:376];
assign DEBUG_select_J_l_GH_BEG1     = ConfigBits[379:378];
assign DEBUG_select_J_l_GH_BEG2     = ConfigBits[381:380];
assign DEBUG_select_J_l_GH_BEG3     = ConfigBits[383:382];
endmodule